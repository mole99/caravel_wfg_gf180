magic
tech gf180mcuC
magscale 1 10
timestamp 1670096641
<< metal1 >>
rect 1344 36874 148624 36908
rect 1344 36822 19624 36874
rect 19676 36822 19728 36874
rect 19780 36822 19832 36874
rect 19884 36822 56444 36874
rect 56496 36822 56548 36874
rect 56600 36822 56652 36874
rect 56704 36822 93264 36874
rect 93316 36822 93368 36874
rect 93420 36822 93472 36874
rect 93524 36822 130084 36874
rect 130136 36822 130188 36874
rect 130240 36822 130292 36874
rect 130344 36822 148624 36874
rect 1344 36788 148624 36822
rect 144162 36542 144174 36594
rect 144226 36542 144238 36594
rect 147746 36542 147758 36594
rect 147810 36542 147822 36594
rect 143042 36430 143054 36482
rect 143106 36430 143118 36482
rect 144834 36430 144846 36482
rect 144898 36430 144910 36482
rect 147074 36430 147086 36482
rect 147138 36430 147150 36482
rect 145954 36318 145966 36370
rect 146018 36318 146030 36370
rect 142158 36258 142210 36270
rect 142158 36194 142210 36206
rect 1344 36090 148784 36124
rect 1344 36038 38034 36090
rect 38086 36038 38138 36090
rect 38190 36038 38242 36090
rect 38294 36038 74854 36090
rect 74906 36038 74958 36090
rect 75010 36038 75062 36090
rect 75114 36038 111674 36090
rect 111726 36038 111778 36090
rect 111830 36038 111882 36090
rect 111934 36038 148494 36090
rect 148546 36038 148598 36090
rect 148650 36038 148702 36090
rect 148754 36038 148784 36090
rect 1344 36004 148784 36038
rect 144946 35646 144958 35698
rect 145010 35646 145022 35698
rect 146738 35646 146750 35698
rect 146802 35646 146814 35698
rect 143838 35586 143890 35598
rect 143838 35522 143890 35534
rect 144286 35586 144338 35598
rect 146066 35534 146078 35586
rect 146130 35534 146142 35586
rect 147634 35534 147646 35586
rect 147698 35534 147710 35586
rect 144286 35522 144338 35534
rect 1344 35306 148624 35340
rect 1344 35254 19624 35306
rect 19676 35254 19728 35306
rect 19780 35254 19832 35306
rect 19884 35254 56444 35306
rect 56496 35254 56548 35306
rect 56600 35254 56652 35306
rect 56704 35254 93264 35306
rect 93316 35254 93368 35306
rect 93420 35254 93472 35306
rect 93524 35254 130084 35306
rect 130136 35254 130188 35306
rect 130240 35254 130292 35306
rect 130344 35254 148624 35306
rect 1344 35220 148624 35254
rect 144946 34862 144958 34914
rect 145010 34862 145022 34914
rect 146066 34750 146078 34802
rect 146130 34750 146142 34802
rect 144398 34690 144450 34702
rect 144398 34626 144450 34638
rect 146638 34690 146690 34702
rect 146638 34626 146690 34638
rect 147086 34690 147138 34702
rect 147086 34626 147138 34638
rect 1344 34522 148784 34556
rect 1344 34470 38034 34522
rect 38086 34470 38138 34522
rect 38190 34470 38242 34522
rect 38294 34470 74854 34522
rect 74906 34470 74958 34522
rect 75010 34470 75062 34522
rect 75114 34470 111674 34522
rect 111726 34470 111778 34522
rect 111830 34470 111882 34522
rect 111934 34470 148494 34522
rect 148546 34470 148598 34522
rect 148650 34470 148702 34522
rect 148754 34470 148784 34522
rect 1344 34436 148784 34470
rect 144946 34078 144958 34130
rect 145010 34078 145022 34130
rect 144286 34018 144338 34030
rect 146066 33966 146078 34018
rect 146130 33966 146142 34018
rect 144286 33954 144338 33966
rect 1344 33738 148624 33772
rect 1344 33686 19624 33738
rect 19676 33686 19728 33738
rect 19780 33686 19832 33738
rect 19884 33686 56444 33738
rect 56496 33686 56548 33738
rect 56600 33686 56652 33738
rect 56704 33686 93264 33738
rect 93316 33686 93368 33738
rect 93420 33686 93472 33738
rect 93524 33686 130084 33738
rect 130136 33686 130188 33738
rect 130240 33686 130292 33738
rect 130344 33686 148624 33738
rect 1344 33652 148624 33686
rect 144946 33294 144958 33346
rect 145010 33294 145022 33346
rect 146066 33182 146078 33234
rect 146130 33182 146142 33234
rect 144398 33122 144450 33134
rect 144398 33058 144450 33070
rect 1344 32954 148784 32988
rect 1344 32902 38034 32954
rect 38086 32902 38138 32954
rect 38190 32902 38242 32954
rect 38294 32902 74854 32954
rect 74906 32902 74958 32954
rect 75010 32902 75062 32954
rect 75114 32902 111674 32954
rect 111726 32902 111778 32954
rect 111830 32902 111882 32954
rect 111934 32902 148494 32954
rect 148546 32902 148598 32954
rect 148650 32902 148702 32954
rect 148754 32902 148784 32954
rect 1344 32868 148784 32902
rect 1344 32170 148624 32204
rect 1344 32118 19624 32170
rect 19676 32118 19728 32170
rect 19780 32118 19832 32170
rect 19884 32118 56444 32170
rect 56496 32118 56548 32170
rect 56600 32118 56652 32170
rect 56704 32118 93264 32170
rect 93316 32118 93368 32170
rect 93420 32118 93472 32170
rect 93524 32118 130084 32170
rect 130136 32118 130188 32170
rect 130240 32118 130292 32170
rect 130344 32118 148624 32170
rect 1344 32084 148624 32118
rect 144946 31726 144958 31778
rect 145010 31726 145022 31778
rect 146066 31614 146078 31666
rect 146130 31614 146142 31666
rect 144398 31554 144450 31566
rect 144398 31490 144450 31502
rect 1344 31386 148784 31420
rect 1344 31334 38034 31386
rect 38086 31334 38138 31386
rect 38190 31334 38242 31386
rect 38294 31334 74854 31386
rect 74906 31334 74958 31386
rect 75010 31334 75062 31386
rect 75114 31334 111674 31386
rect 111726 31334 111778 31386
rect 111830 31334 111882 31386
rect 111934 31334 148494 31386
rect 148546 31334 148598 31386
rect 148650 31334 148702 31386
rect 148754 31334 148784 31386
rect 1344 31300 148784 31334
rect 144946 30942 144958 30994
rect 145010 30942 145022 30994
rect 144286 30882 144338 30894
rect 146066 30830 146078 30882
rect 146130 30830 146142 30882
rect 144286 30818 144338 30830
rect 1344 30602 148624 30636
rect 1344 30550 19624 30602
rect 19676 30550 19728 30602
rect 19780 30550 19832 30602
rect 19884 30550 56444 30602
rect 56496 30550 56548 30602
rect 56600 30550 56652 30602
rect 56704 30550 93264 30602
rect 93316 30550 93368 30602
rect 93420 30550 93472 30602
rect 93524 30550 130084 30602
rect 130136 30550 130188 30602
rect 130240 30550 130292 30602
rect 130344 30550 148624 30602
rect 1344 30516 148624 30550
rect 144946 30158 144958 30210
rect 145010 30158 145022 30210
rect 146066 30046 146078 30098
rect 146130 30046 146142 30098
rect 144398 29986 144450 29998
rect 144398 29922 144450 29934
rect 1344 29818 148784 29852
rect 1344 29766 38034 29818
rect 38086 29766 38138 29818
rect 38190 29766 38242 29818
rect 38294 29766 74854 29818
rect 74906 29766 74958 29818
rect 75010 29766 75062 29818
rect 75114 29766 111674 29818
rect 111726 29766 111778 29818
rect 111830 29766 111882 29818
rect 111934 29766 148494 29818
rect 148546 29766 148598 29818
rect 148650 29766 148702 29818
rect 148754 29766 148784 29818
rect 1344 29732 148784 29766
rect 144946 29374 144958 29426
rect 145010 29374 145022 29426
rect 144286 29314 144338 29326
rect 146066 29262 146078 29314
rect 146130 29262 146142 29314
rect 144286 29250 144338 29262
rect 1344 29034 148624 29068
rect 1344 28982 19624 29034
rect 19676 28982 19728 29034
rect 19780 28982 19832 29034
rect 19884 28982 56444 29034
rect 56496 28982 56548 29034
rect 56600 28982 56652 29034
rect 56704 28982 93264 29034
rect 93316 28982 93368 29034
rect 93420 28982 93472 29034
rect 93524 28982 130084 29034
rect 130136 28982 130188 29034
rect 130240 28982 130292 29034
rect 130344 28982 148624 29034
rect 1344 28948 148624 28982
rect 144398 28642 144450 28654
rect 146078 28642 146130 28654
rect 144946 28590 144958 28642
rect 145010 28590 145022 28642
rect 144398 28578 144450 28590
rect 146078 28578 146130 28590
rect 1344 28250 148784 28284
rect 1344 28198 38034 28250
rect 38086 28198 38138 28250
rect 38190 28198 38242 28250
rect 38294 28198 74854 28250
rect 74906 28198 74958 28250
rect 75010 28198 75062 28250
rect 75114 28198 111674 28250
rect 111726 28198 111778 28250
rect 111830 28198 111882 28250
rect 111934 28198 148494 28250
rect 148546 28198 148598 28250
rect 148650 28198 148702 28250
rect 148754 28198 148784 28250
rect 1344 28164 148784 28198
rect 144946 27806 144958 27858
rect 145010 27806 145022 27858
rect 144286 27746 144338 27758
rect 146066 27694 146078 27746
rect 146130 27694 146142 27746
rect 144286 27682 144338 27694
rect 1344 27466 148624 27500
rect 1344 27414 19624 27466
rect 19676 27414 19728 27466
rect 19780 27414 19832 27466
rect 19884 27414 56444 27466
rect 56496 27414 56548 27466
rect 56600 27414 56652 27466
rect 56704 27414 93264 27466
rect 93316 27414 93368 27466
rect 93420 27414 93472 27466
rect 93524 27414 130084 27466
rect 130136 27414 130188 27466
rect 130240 27414 130292 27466
rect 130344 27414 148624 27466
rect 1344 27380 148624 27414
rect 144946 27022 144958 27074
rect 145010 27022 145022 27074
rect 144398 26962 144450 26974
rect 146066 26910 146078 26962
rect 146130 26910 146142 26962
rect 144398 26898 144450 26910
rect 1344 26682 148784 26716
rect 1344 26630 38034 26682
rect 38086 26630 38138 26682
rect 38190 26630 38242 26682
rect 38294 26630 74854 26682
rect 74906 26630 74958 26682
rect 75010 26630 75062 26682
rect 75114 26630 111674 26682
rect 111726 26630 111778 26682
rect 111830 26630 111882 26682
rect 111934 26630 148494 26682
rect 148546 26630 148598 26682
rect 148650 26630 148702 26682
rect 148754 26630 148784 26682
rect 1344 26596 148784 26630
rect 1344 25898 148624 25932
rect 1344 25846 19624 25898
rect 19676 25846 19728 25898
rect 19780 25846 19832 25898
rect 19884 25846 56444 25898
rect 56496 25846 56548 25898
rect 56600 25846 56652 25898
rect 56704 25846 93264 25898
rect 93316 25846 93368 25898
rect 93420 25846 93472 25898
rect 93524 25846 130084 25898
rect 130136 25846 130188 25898
rect 130240 25846 130292 25898
rect 130344 25846 148624 25898
rect 1344 25812 148624 25846
rect 144946 25454 144958 25506
rect 145010 25454 145022 25506
rect 146066 25342 146078 25394
rect 146130 25342 146142 25394
rect 144398 25282 144450 25294
rect 144398 25218 144450 25230
rect 1344 25114 148784 25148
rect 1344 25062 38034 25114
rect 38086 25062 38138 25114
rect 38190 25062 38242 25114
rect 38294 25062 74854 25114
rect 74906 25062 74958 25114
rect 75010 25062 75062 25114
rect 75114 25062 111674 25114
rect 111726 25062 111778 25114
rect 111830 25062 111882 25114
rect 111934 25062 148494 25114
rect 148546 25062 148598 25114
rect 148650 25062 148702 25114
rect 148754 25062 148784 25114
rect 1344 25028 148784 25062
rect 144946 24670 144958 24722
rect 145010 24670 145022 24722
rect 144286 24610 144338 24622
rect 146066 24558 146078 24610
rect 146130 24558 146142 24610
rect 144286 24546 144338 24558
rect 1344 24330 148624 24364
rect 1344 24278 19624 24330
rect 19676 24278 19728 24330
rect 19780 24278 19832 24330
rect 19884 24278 56444 24330
rect 56496 24278 56548 24330
rect 56600 24278 56652 24330
rect 56704 24278 93264 24330
rect 93316 24278 93368 24330
rect 93420 24278 93472 24330
rect 93524 24278 130084 24330
rect 130136 24278 130188 24330
rect 130240 24278 130292 24330
rect 130344 24278 148624 24330
rect 1344 24244 148624 24278
rect 144946 23886 144958 23938
rect 145010 23886 145022 23938
rect 146066 23774 146078 23826
rect 146130 23774 146142 23826
rect 144398 23714 144450 23726
rect 144398 23650 144450 23662
rect 1344 23546 148784 23580
rect 1344 23494 38034 23546
rect 38086 23494 38138 23546
rect 38190 23494 38242 23546
rect 38294 23494 74854 23546
rect 74906 23494 74958 23546
rect 75010 23494 75062 23546
rect 75114 23494 111674 23546
rect 111726 23494 111778 23546
rect 111830 23494 111882 23546
rect 111934 23494 148494 23546
rect 148546 23494 148598 23546
rect 148650 23494 148702 23546
rect 148754 23494 148784 23546
rect 1344 23460 148784 23494
rect 144946 23102 144958 23154
rect 145010 23102 145022 23154
rect 144286 23042 144338 23054
rect 146066 22990 146078 23042
rect 146130 22990 146142 23042
rect 144286 22978 144338 22990
rect 1344 22762 148624 22796
rect 1344 22710 19624 22762
rect 19676 22710 19728 22762
rect 19780 22710 19832 22762
rect 19884 22710 56444 22762
rect 56496 22710 56548 22762
rect 56600 22710 56652 22762
rect 56704 22710 93264 22762
rect 93316 22710 93368 22762
rect 93420 22710 93472 22762
rect 93524 22710 130084 22762
rect 130136 22710 130188 22762
rect 130240 22710 130292 22762
rect 130344 22710 148624 22762
rect 1344 22676 148624 22710
rect 144946 22318 144958 22370
rect 145010 22318 145022 22370
rect 146066 22206 146078 22258
rect 146130 22206 146142 22258
rect 144398 22146 144450 22158
rect 144398 22082 144450 22094
rect 1344 21978 148784 22012
rect 1344 21926 38034 21978
rect 38086 21926 38138 21978
rect 38190 21926 38242 21978
rect 38294 21926 74854 21978
rect 74906 21926 74958 21978
rect 75010 21926 75062 21978
rect 75114 21926 111674 21978
rect 111726 21926 111778 21978
rect 111830 21926 111882 21978
rect 111934 21926 148494 21978
rect 148546 21926 148598 21978
rect 148650 21926 148702 21978
rect 148754 21926 148784 21978
rect 1344 21892 148784 21926
rect 144946 21534 144958 21586
rect 145010 21534 145022 21586
rect 144286 21474 144338 21486
rect 146066 21422 146078 21474
rect 146130 21422 146142 21474
rect 144286 21410 144338 21422
rect 1344 21194 148624 21228
rect 1344 21142 19624 21194
rect 19676 21142 19728 21194
rect 19780 21142 19832 21194
rect 19884 21142 56444 21194
rect 56496 21142 56548 21194
rect 56600 21142 56652 21194
rect 56704 21142 93264 21194
rect 93316 21142 93368 21194
rect 93420 21142 93472 21194
rect 93524 21142 130084 21194
rect 130136 21142 130188 21194
rect 130240 21142 130292 21194
rect 130344 21142 148624 21194
rect 1344 21108 148624 21142
rect 144946 20750 144958 20802
rect 145010 20750 145022 20802
rect 146066 20638 146078 20690
rect 146130 20638 146142 20690
rect 144398 20578 144450 20590
rect 144398 20514 144450 20526
rect 1344 20410 148784 20444
rect 1344 20358 38034 20410
rect 38086 20358 38138 20410
rect 38190 20358 38242 20410
rect 38294 20358 74854 20410
rect 74906 20358 74958 20410
rect 75010 20358 75062 20410
rect 75114 20358 111674 20410
rect 111726 20358 111778 20410
rect 111830 20358 111882 20410
rect 111934 20358 148494 20410
rect 148546 20358 148598 20410
rect 148650 20358 148702 20410
rect 148754 20358 148784 20410
rect 1344 20324 148784 20358
rect 1344 19626 148624 19660
rect 1344 19574 19624 19626
rect 19676 19574 19728 19626
rect 19780 19574 19832 19626
rect 19884 19574 56444 19626
rect 56496 19574 56548 19626
rect 56600 19574 56652 19626
rect 56704 19574 93264 19626
rect 93316 19574 93368 19626
rect 93420 19574 93472 19626
rect 93524 19574 130084 19626
rect 130136 19574 130188 19626
rect 130240 19574 130292 19626
rect 130344 19574 148624 19626
rect 1344 19540 148624 19574
rect 144946 19182 144958 19234
rect 145010 19182 145022 19234
rect 146066 19070 146078 19122
rect 146130 19070 146142 19122
rect 144398 19010 144450 19022
rect 144398 18946 144450 18958
rect 1344 18842 148784 18876
rect 1344 18790 38034 18842
rect 38086 18790 38138 18842
rect 38190 18790 38242 18842
rect 38294 18790 74854 18842
rect 74906 18790 74958 18842
rect 75010 18790 75062 18842
rect 75114 18790 111674 18842
rect 111726 18790 111778 18842
rect 111830 18790 111882 18842
rect 111934 18790 148494 18842
rect 148546 18790 148598 18842
rect 148650 18790 148702 18842
rect 148754 18790 148784 18842
rect 1344 18756 148784 18790
rect 111582 18674 111634 18686
rect 111582 18610 111634 18622
rect 111246 18562 111298 18574
rect 111246 18498 111298 18510
rect 144946 18398 144958 18450
rect 145010 18398 145022 18450
rect 110686 18338 110738 18350
rect 110686 18274 110738 18286
rect 144286 18338 144338 18350
rect 146066 18286 146078 18338
rect 146130 18286 146142 18338
rect 144286 18274 144338 18286
rect 1344 18058 148624 18092
rect 1344 18006 19624 18058
rect 19676 18006 19728 18058
rect 19780 18006 19832 18058
rect 19884 18006 56444 18058
rect 56496 18006 56548 18058
rect 56600 18006 56652 18058
rect 56704 18006 93264 18058
rect 93316 18006 93368 18058
rect 93420 18006 93472 18058
rect 93524 18006 130084 18058
rect 130136 18006 130188 18058
rect 130240 18006 130292 18058
rect 130344 18006 148624 18058
rect 1344 17972 148624 18006
rect 144946 17614 144958 17666
rect 145010 17614 145022 17666
rect 146066 17502 146078 17554
rect 146130 17502 146142 17554
rect 144398 17442 144450 17454
rect 144398 17378 144450 17390
rect 1344 17274 148784 17308
rect 1344 17222 38034 17274
rect 38086 17222 38138 17274
rect 38190 17222 38242 17274
rect 38294 17222 74854 17274
rect 74906 17222 74958 17274
rect 75010 17222 75062 17274
rect 75114 17222 111674 17274
rect 111726 17222 111778 17274
rect 111830 17222 111882 17274
rect 111934 17222 148494 17274
rect 148546 17222 148598 17274
rect 148650 17222 148702 17274
rect 148754 17222 148784 17274
rect 1344 17188 148784 17222
rect 144286 16882 144338 16894
rect 146078 16882 146130 16894
rect 144946 16830 144958 16882
rect 145010 16830 145022 16882
rect 144286 16818 144338 16830
rect 146078 16818 146130 16830
rect 1344 16490 148624 16524
rect 1344 16438 19624 16490
rect 19676 16438 19728 16490
rect 19780 16438 19832 16490
rect 19884 16438 56444 16490
rect 56496 16438 56548 16490
rect 56600 16438 56652 16490
rect 56704 16438 93264 16490
rect 93316 16438 93368 16490
rect 93420 16438 93472 16490
rect 93524 16438 130084 16490
rect 130136 16438 130188 16490
rect 130240 16438 130292 16490
rect 130344 16438 148624 16490
rect 1344 16404 148624 16438
rect 144946 16046 144958 16098
rect 145010 16046 145022 16098
rect 146066 15934 146078 15986
rect 146130 15934 146142 15986
rect 144398 15874 144450 15886
rect 144398 15810 144450 15822
rect 1344 15706 148784 15740
rect 1344 15654 38034 15706
rect 38086 15654 38138 15706
rect 38190 15654 38242 15706
rect 38294 15654 74854 15706
rect 74906 15654 74958 15706
rect 75010 15654 75062 15706
rect 75114 15654 111674 15706
rect 111726 15654 111778 15706
rect 111830 15654 111882 15706
rect 111934 15654 148494 15706
rect 148546 15654 148598 15706
rect 148650 15654 148702 15706
rect 148754 15654 148784 15706
rect 1344 15620 148784 15654
rect 144946 15262 144958 15314
rect 145010 15262 145022 15314
rect 144286 15202 144338 15214
rect 146066 15150 146078 15202
rect 146130 15150 146142 15202
rect 144286 15138 144338 15150
rect 1344 14922 148624 14956
rect 1344 14870 19624 14922
rect 19676 14870 19728 14922
rect 19780 14870 19832 14922
rect 19884 14870 56444 14922
rect 56496 14870 56548 14922
rect 56600 14870 56652 14922
rect 56704 14870 93264 14922
rect 93316 14870 93368 14922
rect 93420 14870 93472 14922
rect 93524 14870 130084 14922
rect 130136 14870 130188 14922
rect 130240 14870 130292 14922
rect 130344 14870 148624 14922
rect 1344 14836 148624 14870
rect 144946 14478 144958 14530
rect 145010 14478 145022 14530
rect 146066 14366 146078 14418
rect 146130 14366 146142 14418
rect 144398 14306 144450 14318
rect 144398 14242 144450 14254
rect 1344 14138 148784 14172
rect 1344 14086 38034 14138
rect 38086 14086 38138 14138
rect 38190 14086 38242 14138
rect 38294 14086 74854 14138
rect 74906 14086 74958 14138
rect 75010 14086 75062 14138
rect 75114 14086 111674 14138
rect 111726 14086 111778 14138
rect 111830 14086 111882 14138
rect 111934 14086 148494 14138
rect 148546 14086 148598 14138
rect 148650 14086 148702 14138
rect 148754 14086 148784 14138
rect 1344 14052 148784 14086
rect 1344 13354 148624 13388
rect 1344 13302 19624 13354
rect 19676 13302 19728 13354
rect 19780 13302 19832 13354
rect 19884 13302 56444 13354
rect 56496 13302 56548 13354
rect 56600 13302 56652 13354
rect 56704 13302 93264 13354
rect 93316 13302 93368 13354
rect 93420 13302 93472 13354
rect 93524 13302 130084 13354
rect 130136 13302 130188 13354
rect 130240 13302 130292 13354
rect 130344 13302 148624 13354
rect 1344 13268 148624 13302
rect 144946 12910 144958 12962
rect 145010 12910 145022 12962
rect 101166 12850 101218 12862
rect 101166 12786 101218 12798
rect 101502 12850 101554 12862
rect 146066 12798 146078 12850
rect 146130 12798 146142 12850
rect 101502 12786 101554 12798
rect 144398 12738 144450 12750
rect 144398 12674 144450 12686
rect 1344 12570 148784 12604
rect 1344 12518 38034 12570
rect 38086 12518 38138 12570
rect 38190 12518 38242 12570
rect 38294 12518 74854 12570
rect 74906 12518 74958 12570
rect 75010 12518 75062 12570
rect 75114 12518 111674 12570
rect 111726 12518 111778 12570
rect 111830 12518 111882 12570
rect 111934 12518 148494 12570
rect 148546 12518 148598 12570
rect 148650 12518 148702 12570
rect 148754 12518 148784 12570
rect 1344 12484 148784 12518
rect 100494 12402 100546 12414
rect 100494 12338 100546 12350
rect 100158 12178 100210 12190
rect 144946 12126 144958 12178
rect 145010 12126 145022 12178
rect 100158 12114 100210 12126
rect 144286 12066 144338 12078
rect 146066 12014 146078 12066
rect 146130 12014 146142 12066
rect 144286 12002 144338 12014
rect 1344 11786 148624 11820
rect 1344 11734 19624 11786
rect 19676 11734 19728 11786
rect 19780 11734 19832 11786
rect 19884 11734 56444 11786
rect 56496 11734 56548 11786
rect 56600 11734 56652 11786
rect 56704 11734 93264 11786
rect 93316 11734 93368 11786
rect 93420 11734 93472 11786
rect 93524 11734 130084 11786
rect 130136 11734 130188 11786
rect 130240 11734 130292 11786
rect 130344 11734 148624 11786
rect 1344 11700 148624 11734
rect 144946 11342 144958 11394
rect 145010 11342 145022 11394
rect 101166 11282 101218 11294
rect 146066 11230 146078 11282
rect 146130 11230 146142 11282
rect 101166 11218 101218 11230
rect 100494 11170 100546 11182
rect 100494 11106 100546 11118
rect 101502 11170 101554 11182
rect 101502 11106 101554 11118
rect 144398 11170 144450 11182
rect 144398 11106 144450 11118
rect 1344 11002 148784 11036
rect 1344 10950 38034 11002
rect 38086 10950 38138 11002
rect 38190 10950 38242 11002
rect 38294 10950 74854 11002
rect 74906 10950 74958 11002
rect 75010 10950 75062 11002
rect 75114 10950 111674 11002
rect 111726 10950 111778 11002
rect 111830 10950 111882 11002
rect 111934 10950 148494 11002
rect 148546 10950 148598 11002
rect 148650 10950 148702 11002
rect 148754 10950 148784 11002
rect 1344 10916 148784 10950
rect 146290 10670 146302 10722
rect 146354 10670 146366 10722
rect 146862 10498 146914 10510
rect 145170 10446 145182 10498
rect 145234 10446 145246 10498
rect 146862 10434 146914 10446
rect 1344 10218 148624 10252
rect 1344 10166 19624 10218
rect 19676 10166 19728 10218
rect 19780 10166 19832 10218
rect 19884 10166 56444 10218
rect 56496 10166 56548 10218
rect 56600 10166 56652 10218
rect 56704 10166 93264 10218
rect 93316 10166 93368 10218
rect 93420 10166 93472 10218
rect 93524 10166 130084 10218
rect 130136 10166 130188 10218
rect 130240 10166 130292 10218
rect 130344 10166 148624 10218
rect 1344 10132 148624 10166
rect 144946 9886 144958 9938
rect 145010 9886 145022 9938
rect 146290 9662 146302 9714
rect 146354 9662 146366 9714
rect 146974 9602 147026 9614
rect 146974 9538 147026 9550
rect 1344 9434 148784 9468
rect 1344 9382 38034 9434
rect 38086 9382 38138 9434
rect 38190 9382 38242 9434
rect 38294 9382 74854 9434
rect 74906 9382 74958 9434
rect 75010 9382 75062 9434
rect 75114 9382 111674 9434
rect 111726 9382 111778 9434
rect 111830 9382 111882 9434
rect 111934 9382 148494 9434
rect 148546 9382 148598 9434
rect 148650 9382 148702 9434
rect 148754 9382 148784 9434
rect 1344 9348 148784 9382
rect 146290 9102 146302 9154
rect 146354 9102 146366 9154
rect 146862 8930 146914 8942
rect 144946 8878 144958 8930
rect 145010 8878 145022 8930
rect 146862 8866 146914 8878
rect 1344 8650 148624 8684
rect 1344 8598 19624 8650
rect 19676 8598 19728 8650
rect 19780 8598 19832 8650
rect 19884 8598 56444 8650
rect 56496 8598 56548 8650
rect 56600 8598 56652 8650
rect 56704 8598 93264 8650
rect 93316 8598 93368 8650
rect 93420 8598 93472 8650
rect 93524 8598 130084 8650
rect 130136 8598 130188 8650
rect 130240 8598 130292 8650
rect 130344 8598 148624 8650
rect 1344 8564 148624 8598
rect 144946 8318 144958 8370
rect 145010 8318 145022 8370
rect 146290 8094 146302 8146
rect 146354 8094 146366 8146
rect 146974 8034 147026 8046
rect 146974 7970 147026 7982
rect 1344 7866 148784 7900
rect 1344 7814 38034 7866
rect 38086 7814 38138 7866
rect 38190 7814 38242 7866
rect 38294 7814 74854 7866
rect 74906 7814 74958 7866
rect 75010 7814 75062 7866
rect 75114 7814 111674 7866
rect 111726 7814 111778 7866
rect 111830 7814 111882 7866
rect 111934 7814 148494 7866
rect 148546 7814 148598 7866
rect 148650 7814 148702 7866
rect 148754 7814 148784 7866
rect 1344 7780 148784 7814
rect 105534 7698 105586 7710
rect 105534 7634 105586 7646
rect 139022 7698 139074 7710
rect 139022 7634 139074 7646
rect 139918 7698 139970 7710
rect 139918 7634 139970 7646
rect 129838 7586 129890 7598
rect 129838 7522 129890 7534
rect 130958 7586 131010 7598
rect 130958 7522 131010 7534
rect 131294 7586 131346 7598
rect 131294 7522 131346 7534
rect 131742 7586 131794 7598
rect 146862 7586 146914 7598
rect 146178 7534 146190 7586
rect 146242 7534 146254 7586
rect 131742 7522 131794 7534
rect 146862 7522 146914 7534
rect 105298 7422 105310 7474
rect 105362 7422 105374 7474
rect 138786 7422 138798 7474
rect 138850 7422 138862 7474
rect 139682 7422 139694 7474
rect 139746 7422 139758 7474
rect 130398 7362 130450 7374
rect 130398 7298 130450 7310
rect 137790 7362 137842 7374
rect 137790 7298 137842 7310
rect 140366 7362 140418 7374
rect 140366 7298 140418 7310
rect 144286 7362 144338 7374
rect 144946 7310 144958 7362
rect 145010 7310 145022 7362
rect 144286 7298 144338 7310
rect 130386 7198 130398 7250
rect 130450 7247 130462 7250
rect 130610 7247 130622 7250
rect 130450 7201 130622 7247
rect 130450 7198 130462 7201
rect 130610 7198 130622 7201
rect 130674 7198 130686 7250
rect 1344 7082 148624 7116
rect 1344 7030 19624 7082
rect 19676 7030 19728 7082
rect 19780 7030 19832 7082
rect 19884 7030 56444 7082
rect 56496 7030 56548 7082
rect 56600 7030 56652 7082
rect 56704 7030 93264 7082
rect 93316 7030 93368 7082
rect 93420 7030 93472 7082
rect 93524 7030 130084 7082
rect 130136 7030 130188 7082
rect 130240 7030 130292 7082
rect 130344 7030 148624 7082
rect 1344 6996 148624 7030
rect 139246 6914 139298 6926
rect 139246 6850 139298 6862
rect 138910 6802 138962 6814
rect 142930 6750 142942 6802
rect 142994 6750 143006 6802
rect 145058 6750 145070 6802
rect 145122 6750 145134 6802
rect 138910 6738 138962 6750
rect 110462 6690 110514 6702
rect 110462 6626 110514 6638
rect 117966 6690 118018 6702
rect 117966 6626 118018 6638
rect 128830 6690 128882 6702
rect 128830 6626 128882 6638
rect 129614 6690 129666 6702
rect 129614 6626 129666 6638
rect 131966 6690 132018 6702
rect 131966 6626 132018 6638
rect 137566 6690 137618 6702
rect 137566 6626 137618 6638
rect 139918 6690 139970 6702
rect 139918 6626 139970 6638
rect 101166 6578 101218 6590
rect 101166 6514 101218 6526
rect 101502 6578 101554 6590
rect 101502 6514 101554 6526
rect 103294 6578 103346 6590
rect 103294 6514 103346 6526
rect 103630 6578 103682 6590
rect 103630 6514 103682 6526
rect 104190 6578 104242 6590
rect 104190 6514 104242 6526
rect 104526 6578 104578 6590
rect 104526 6514 104578 6526
rect 105198 6578 105250 6590
rect 105198 6514 105250 6526
rect 105534 6578 105586 6590
rect 105534 6514 105586 6526
rect 117070 6578 117122 6590
rect 117070 6514 117122 6526
rect 117406 6578 117458 6590
rect 117406 6514 117458 6526
rect 130174 6578 130226 6590
rect 130174 6514 130226 6526
rect 130510 6578 130562 6590
rect 130510 6514 130562 6526
rect 131070 6578 131122 6590
rect 131070 6514 131122 6526
rect 131406 6578 131458 6590
rect 131406 6514 131458 6526
rect 132974 6578 133026 6590
rect 132974 6514 133026 6526
rect 133310 6578 133362 6590
rect 140926 6578 140978 6590
rect 138114 6526 138126 6578
rect 138178 6526 138190 6578
rect 138674 6526 138686 6578
rect 138738 6526 138750 6578
rect 133310 6514 133362 6526
rect 140926 6514 140978 6526
rect 141262 6578 141314 6590
rect 146974 6578 147026 6590
rect 144274 6526 144286 6578
rect 144338 6526 144350 6578
rect 146290 6526 146302 6578
rect 146354 6526 146366 6578
rect 141262 6514 141314 6526
rect 146974 6514 147026 6526
rect 105982 6466 106034 6478
rect 105982 6402 106034 6414
rect 111022 6466 111074 6478
rect 111022 6402 111074 6414
rect 111470 6466 111522 6478
rect 111470 6402 111522 6414
rect 112702 6466 112754 6478
rect 112702 6402 112754 6414
rect 124350 6466 124402 6478
rect 124350 6402 124402 6414
rect 129278 6466 129330 6478
rect 129278 6402 129330 6414
rect 133982 6466 134034 6478
rect 133982 6402 134034 6414
rect 137006 6466 137058 6478
rect 137006 6402 137058 6414
rect 1344 6298 148784 6332
rect 1344 6246 38034 6298
rect 38086 6246 38138 6298
rect 38190 6246 38242 6298
rect 38294 6246 74854 6298
rect 74906 6246 74958 6298
rect 75010 6246 75062 6298
rect 75114 6246 111674 6298
rect 111726 6246 111778 6298
rect 111830 6246 111882 6298
rect 111934 6246 148494 6298
rect 148546 6246 148598 6298
rect 148650 6246 148702 6298
rect 148754 6246 148784 6298
rect 1344 6212 148784 6246
rect 82798 6130 82850 6142
rect 82798 6066 82850 6078
rect 86942 6130 86994 6142
rect 86942 6066 86994 6078
rect 88398 6130 88450 6142
rect 88398 6066 88450 6078
rect 98478 6130 98530 6142
rect 98478 6066 98530 6078
rect 101950 6130 102002 6142
rect 101950 6066 102002 6078
rect 103742 6130 103794 6142
rect 103742 6066 103794 6078
rect 105310 6130 105362 6142
rect 105310 6066 105362 6078
rect 106990 6130 107042 6142
rect 106990 6066 107042 6078
rect 109118 6130 109170 6142
rect 109118 6066 109170 6078
rect 110910 6130 110962 6142
rect 110910 6066 110962 6078
rect 113486 6130 113538 6142
rect 113486 6066 113538 6078
rect 115278 6130 115330 6142
rect 115278 6066 115330 6078
rect 120094 6130 120146 6142
rect 120094 6066 120146 6078
rect 122110 6130 122162 6142
rect 122110 6066 122162 6078
rect 124910 6130 124962 6142
rect 124910 6066 124962 6078
rect 126030 6130 126082 6142
rect 126030 6066 126082 6078
rect 130510 6130 130562 6142
rect 130510 6066 130562 6078
rect 134766 6130 134818 6142
rect 134766 6066 134818 6078
rect 136222 6130 136274 6142
rect 136222 6066 136274 6078
rect 137342 6130 137394 6142
rect 137342 6066 137394 6078
rect 141150 6130 141202 6142
rect 141150 6066 141202 6078
rect 142158 6130 142210 6142
rect 142158 6066 142210 6078
rect 112030 6018 112082 6030
rect 97458 5966 97470 6018
rect 97522 5966 97534 6018
rect 97906 5966 97918 6018
rect 97970 5966 97982 6018
rect 102722 5966 102734 6018
rect 102786 5966 102798 6018
rect 106194 5966 106206 6018
rect 106258 5966 106270 6018
rect 109890 5966 109902 6018
rect 109954 5966 109966 6018
rect 116050 5966 116062 6018
rect 116114 5966 116126 6018
rect 116498 5966 116510 6018
rect 116562 5966 116574 6018
rect 118066 5966 118078 6018
rect 118130 5966 118142 6018
rect 122882 5966 122894 6018
rect 122946 5966 122958 6018
rect 123330 5966 123342 6018
rect 123394 5966 123406 6018
rect 129490 5966 129502 6018
rect 129554 5966 129566 6018
rect 129938 5966 129950 6018
rect 130002 5966 130014 6018
rect 131730 5966 131742 6018
rect 131794 5966 131806 6018
rect 132066 5966 132078 6018
rect 132130 5966 132142 6018
rect 138226 5966 138238 6018
rect 138290 5966 138302 6018
rect 138674 5966 138686 6018
rect 138738 5966 138750 6018
rect 140130 5966 140142 6018
rect 140194 5966 140206 6018
rect 144050 5966 144062 6018
rect 144114 5966 144126 6018
rect 146290 5966 146302 6018
rect 146354 5966 146366 6018
rect 112030 5954 112082 5966
rect 119086 5906 119138 5918
rect 102610 5854 102622 5906
rect 102674 5854 102686 5906
rect 106418 5854 106430 5906
rect 106482 5854 106494 5906
rect 109778 5854 109790 5906
rect 109842 5854 109854 5906
rect 111794 5854 111806 5906
rect 111858 5854 111870 5906
rect 113250 5854 113262 5906
rect 113314 5854 113326 5906
rect 117954 5854 117966 5906
rect 118018 5854 118030 5906
rect 119086 5842 119138 5854
rect 119758 5906 119810 5918
rect 119758 5842 119810 5854
rect 123902 5906 123954 5918
rect 123902 5842 123954 5854
rect 124574 5906 124626 5918
rect 132638 5906 132690 5918
rect 125794 5854 125806 5906
rect 125858 5854 125870 5906
rect 124574 5842 124626 5854
rect 132638 5842 132690 5854
rect 133310 5906 133362 5918
rect 133310 5842 133362 5854
rect 134430 5906 134482 5918
rect 134430 5842 134482 5854
rect 137006 5906 137058 5918
rect 141822 5906 141874 5918
rect 140354 5854 140366 5906
rect 140418 5854 140430 5906
rect 137006 5842 137058 5854
rect 141822 5842 141874 5854
rect 75742 5794 75794 5806
rect 75742 5730 75794 5742
rect 86046 5794 86098 5806
rect 86046 5730 86098 5742
rect 96462 5794 96514 5806
rect 96462 5730 96514 5742
rect 99038 5794 99090 5806
rect 99038 5730 99090 5742
rect 99486 5794 99538 5806
rect 99486 5730 99538 5742
rect 101502 5794 101554 5806
rect 101502 5730 101554 5742
rect 104414 5794 104466 5806
rect 104414 5730 104466 5742
rect 107438 5794 107490 5806
rect 107438 5730 107490 5742
rect 107886 5794 107938 5806
rect 107886 5730 107938 5742
rect 108782 5794 108834 5806
rect 108782 5730 108834 5742
rect 114718 5794 114770 5806
rect 114718 5730 114770 5742
rect 126590 5794 126642 5806
rect 126590 5730 126642 5742
rect 127822 5794 127874 5806
rect 127822 5730 127874 5742
rect 128270 5794 128322 5806
rect 135886 5794 135938 5806
rect 146862 5794 146914 5806
rect 133746 5742 133758 5794
rect 133810 5742 133822 5794
rect 142706 5742 142718 5794
rect 142770 5742 142782 5794
rect 144946 5742 144958 5794
rect 145010 5742 145022 5794
rect 128270 5730 128322 5742
rect 135886 5730 135938 5742
rect 146862 5730 146914 5742
rect 147310 5794 147362 5806
rect 147310 5730 147362 5742
rect 98142 5682 98194 5694
rect 98142 5618 98194 5630
rect 103406 5682 103458 5694
rect 103406 5618 103458 5630
rect 105646 5682 105698 5694
rect 110574 5682 110626 5694
rect 106754 5630 106766 5682
rect 106818 5679 106830 5682
rect 107426 5679 107438 5682
rect 106818 5633 107438 5679
rect 106818 5630 106830 5633
rect 107426 5630 107438 5633
rect 107490 5630 107502 5682
rect 105646 5618 105698 5630
rect 110574 5618 110626 5630
rect 116734 5682 116786 5694
rect 116734 5618 116786 5630
rect 117070 5682 117122 5694
rect 117070 5618 117122 5630
rect 118750 5682 118802 5694
rect 118750 5618 118802 5630
rect 123566 5682 123618 5694
rect 123566 5618 123618 5630
rect 130174 5682 130226 5694
rect 130174 5618 130226 5630
rect 132302 5682 132354 5694
rect 132302 5618 132354 5630
rect 138910 5682 138962 5694
rect 138910 5618 138962 5630
rect 139246 5682 139298 5694
rect 139246 5618 139298 5630
rect 140814 5682 140866 5694
rect 140814 5618 140866 5630
rect 1344 5514 148624 5548
rect 1344 5462 19624 5514
rect 19676 5462 19728 5514
rect 19780 5462 19832 5514
rect 19884 5462 56444 5514
rect 56496 5462 56548 5514
rect 56600 5462 56652 5514
rect 56704 5462 93264 5514
rect 93316 5462 93368 5514
rect 93420 5462 93472 5514
rect 93524 5462 130084 5514
rect 130136 5462 130188 5514
rect 130240 5462 130292 5514
rect 130344 5462 148624 5514
rect 1344 5428 148624 5462
rect 96238 5346 96290 5358
rect 96238 5282 96290 5294
rect 98142 5346 98194 5358
rect 98142 5282 98194 5294
rect 100046 5346 100098 5358
rect 100046 5282 100098 5294
rect 102958 5346 103010 5358
rect 102958 5282 103010 5294
rect 104862 5346 104914 5358
rect 104862 5282 104914 5294
rect 112254 5346 112306 5358
rect 112254 5282 112306 5294
rect 114158 5346 114210 5358
rect 114158 5282 114210 5294
rect 116174 5346 116226 5358
rect 116174 5282 116226 5294
rect 126254 5346 126306 5358
rect 126254 5282 126306 5294
rect 129726 5346 129778 5358
rect 129726 5282 129778 5294
rect 131742 5346 131794 5358
rect 131742 5282 131794 5294
rect 135438 5346 135490 5358
rect 135438 5282 135490 5294
rect 137342 5346 137394 5358
rect 137342 5282 137394 5294
rect 139246 5346 139298 5358
rect 139246 5282 139298 5294
rect 76190 5234 76242 5246
rect 65650 5182 65662 5234
rect 65714 5182 65726 5234
rect 76190 5170 76242 5182
rect 77646 5234 77698 5246
rect 77646 5170 77698 5182
rect 79438 5234 79490 5246
rect 79438 5170 79490 5182
rect 89854 5234 89906 5246
rect 89854 5170 89906 5182
rect 90302 5234 90354 5246
rect 90302 5170 90354 5182
rect 90750 5234 90802 5246
rect 142930 5182 142942 5234
rect 142994 5182 143006 5234
rect 144946 5182 144958 5234
rect 145010 5182 145022 5234
rect 90750 5170 90802 5182
rect 63758 5122 63810 5134
rect 63758 5058 63810 5070
rect 78542 5122 78594 5134
rect 78542 5058 78594 5070
rect 81006 5122 81058 5134
rect 81006 5058 81058 5070
rect 81454 5122 81506 5134
rect 83358 5122 83410 5134
rect 82226 5070 82238 5122
rect 82290 5070 82302 5122
rect 81454 5058 81506 5070
rect 83358 5058 83410 5070
rect 83806 5122 83858 5134
rect 83806 5058 83858 5070
rect 86718 5122 86770 5134
rect 86718 5058 86770 5070
rect 89406 5122 89458 5134
rect 95902 5122 95954 5134
rect 97806 5122 97858 5134
rect 99710 5122 99762 5134
rect 95442 5070 95454 5122
rect 95506 5070 95518 5122
rect 97346 5070 97358 5122
rect 97410 5070 97422 5122
rect 99250 5070 99262 5122
rect 99314 5070 99326 5122
rect 89406 5058 89458 5070
rect 95902 5058 95954 5070
rect 97806 5058 97858 5070
rect 99710 5058 99762 5070
rect 101054 5122 101106 5134
rect 102622 5122 102674 5134
rect 104526 5122 104578 5134
rect 106430 5122 106482 5134
rect 110014 5122 110066 5134
rect 111918 5122 111970 5134
rect 113822 5122 113874 5134
rect 115838 5122 115890 5134
rect 102162 5070 102174 5122
rect 102226 5070 102238 5122
rect 103730 5070 103742 5122
rect 103794 5070 103806 5122
rect 105858 5070 105870 5122
rect 105922 5070 105934 5122
rect 109554 5070 109566 5122
rect 109618 5070 109630 5122
rect 111458 5070 111470 5122
rect 111522 5070 111534 5122
rect 113138 5070 113150 5122
rect 113202 5070 113214 5122
rect 115378 5070 115390 5122
rect 115442 5070 115454 5122
rect 101054 5058 101106 5070
rect 102622 5058 102674 5070
rect 104526 5058 104578 5070
rect 106430 5058 106482 5070
rect 110014 5058 110066 5070
rect 111918 5058 111970 5070
rect 113822 5058 113874 5070
rect 115838 5058 115890 5070
rect 117966 5122 118018 5134
rect 122782 5122 122834 5134
rect 125918 5122 125970 5134
rect 129390 5122 129442 5134
rect 131406 5122 131458 5134
rect 122322 5070 122334 5122
rect 122386 5070 122398 5122
rect 125458 5070 125470 5122
rect 125522 5070 125534 5122
rect 128930 5070 128942 5122
rect 128994 5070 129006 5122
rect 130946 5070 130958 5122
rect 131010 5070 131022 5122
rect 117966 5058 118018 5070
rect 122782 5058 122834 5070
rect 125918 5058 125970 5070
rect 129390 5058 129442 5070
rect 131406 5058 131458 5070
rect 133534 5122 133586 5134
rect 135102 5122 135154 5134
rect 137006 5122 137058 5134
rect 138910 5122 138962 5134
rect 134642 5070 134654 5122
rect 134706 5070 134718 5122
rect 136546 5070 136558 5122
rect 136610 5070 136622 5122
rect 138450 5070 138462 5122
rect 138514 5070 138526 5122
rect 133534 5058 133586 5070
rect 135102 5058 135154 5070
rect 137006 5058 137058 5070
rect 138910 5058 138962 5070
rect 139806 5122 139858 5134
rect 141822 5122 141874 5134
rect 141138 5070 141150 5122
rect 141202 5070 141214 5122
rect 139806 5058 139858 5070
rect 141822 5058 141874 5070
rect 146862 5122 146914 5134
rect 146862 5058 146914 5070
rect 75406 5010 75458 5022
rect 64306 4958 64318 5010
rect 64370 4958 64382 5010
rect 75406 4946 75458 4958
rect 80670 5010 80722 5022
rect 80670 4946 80722 4958
rect 85486 5010 85538 5022
rect 85486 4946 85538 4958
rect 87726 5010 87778 5022
rect 106766 5010 106818 5022
rect 95106 4958 95118 5010
rect 95170 4958 95182 5010
rect 97010 4958 97022 5010
rect 97074 4958 97086 5010
rect 98914 4958 98926 5010
rect 98978 4958 98990 5010
rect 101826 4958 101838 5010
rect 101890 4958 101902 5010
rect 103954 4958 103966 5010
rect 104018 4958 104030 5010
rect 105634 4958 105646 5010
rect 105698 4958 105710 5010
rect 87726 4946 87778 4958
rect 106766 4946 106818 4958
rect 107438 5010 107490 5022
rect 107438 4946 107490 4958
rect 107774 5010 107826 5022
rect 118302 5010 118354 5022
rect 109218 4958 109230 5010
rect 109282 4958 109294 5010
rect 111122 4958 111134 5010
rect 111186 4958 111198 5010
rect 113026 4958 113038 5010
rect 113090 4958 113102 5010
rect 115042 4958 115054 5010
rect 115106 4958 115118 5010
rect 117170 4958 117182 5010
rect 117234 4958 117246 5010
rect 117730 4958 117742 5010
rect 117794 4958 117806 5010
rect 107774 4946 107826 4958
rect 118302 4946 118354 4958
rect 118974 5010 119026 5022
rect 118974 4946 119026 4958
rect 119310 5010 119362 5022
rect 119310 4946 119362 4958
rect 119870 5010 119922 5022
rect 119870 4946 119922 4958
rect 120206 5010 120258 5022
rect 123118 5010 123170 5022
rect 121986 4958 121998 5010
rect 122050 4958 122062 5010
rect 120206 4946 120258 4958
rect 123118 4946 123170 4958
rect 123790 5010 123842 5022
rect 123790 4946 123842 4958
rect 124126 5010 124178 5022
rect 126814 5010 126866 5022
rect 125122 4958 125134 5010
rect 125186 4958 125198 5010
rect 124126 4946 124178 4958
rect 126814 4946 126866 4958
rect 127598 5010 127650 5022
rect 127598 4946 127650 4958
rect 127934 5010 127986 5022
rect 132974 5010 133026 5022
rect 128818 4958 128830 5010
rect 128882 4958 128894 5010
rect 130610 4958 130622 5010
rect 130674 4958 130686 5010
rect 134418 4958 134430 5010
rect 134482 4958 134494 5010
rect 136434 4958 136446 5010
rect 136498 4958 136510 5010
rect 138338 4958 138350 5010
rect 138402 4958 138414 5010
rect 141250 4958 141262 5010
rect 141314 4958 141326 5010
rect 144274 4958 144286 5010
rect 144338 4958 144350 5010
rect 146290 4958 146302 5010
rect 146354 4958 146366 5010
rect 127934 4946 127986 4958
rect 132974 4946 133026 4958
rect 30382 4898 30434 4910
rect 30382 4834 30434 4846
rect 45502 4898 45554 4910
rect 45502 4834 45554 4846
rect 56926 4898 56978 4910
rect 56926 4834 56978 4846
rect 69358 4898 69410 4910
rect 69358 4834 69410 4846
rect 75742 4898 75794 4910
rect 75742 4834 75794 4846
rect 82462 4898 82514 4910
rect 82462 4834 82514 4846
rect 83022 4898 83074 4910
rect 83022 4834 83074 4846
rect 85822 4898 85874 4910
rect 85822 4834 85874 4846
rect 86382 4898 86434 4910
rect 86382 4834 86434 4846
rect 87390 4898 87442 4910
rect 87390 4834 87442 4846
rect 88174 4898 88226 4910
rect 88174 4834 88226 4846
rect 89070 4898 89122 4910
rect 89070 4834 89122 4846
rect 94558 4898 94610 4910
rect 94558 4834 94610 4846
rect 108222 4898 108274 4910
rect 108222 4834 108274 4846
rect 110350 4898 110402 4910
rect 110350 4834 110402 4846
rect 121438 4898 121490 4910
rect 121438 4834 121490 4846
rect 142158 4898 142210 4910
rect 142158 4834 142210 4846
rect 147422 4898 147474 4910
rect 147422 4834 147474 4846
rect 1344 4730 148784 4764
rect 1344 4678 38034 4730
rect 38086 4678 38138 4730
rect 38190 4678 38242 4730
rect 38294 4678 74854 4730
rect 74906 4678 74958 4730
rect 75010 4678 75062 4730
rect 75114 4678 111674 4730
rect 111726 4678 111778 4730
rect 111830 4678 111882 4730
rect 111934 4678 148494 4730
rect 148546 4678 148598 4730
rect 148650 4678 148702 4730
rect 148754 4678 148784 4730
rect 1344 4644 148784 4678
rect 9774 4562 9826 4574
rect 9774 4498 9826 4510
rect 11342 4562 11394 4574
rect 11342 4498 11394 4510
rect 13022 4562 13074 4574
rect 13022 4498 13074 4510
rect 17054 4562 17106 4574
rect 17054 4498 17106 4510
rect 76526 4562 76578 4574
rect 76526 4498 76578 4510
rect 77982 4562 78034 4574
rect 77982 4498 78034 4510
rect 79774 4562 79826 4574
rect 79774 4498 79826 4510
rect 85374 4562 85426 4574
rect 85374 4498 85426 4510
rect 96462 4562 96514 4574
rect 96462 4498 96514 4510
rect 97134 4562 97186 4574
rect 97134 4498 97186 4510
rect 107102 4562 107154 4574
rect 107102 4498 107154 4510
rect 120206 4562 120258 4574
rect 120206 4498 120258 4510
rect 123454 4562 123506 4574
rect 123454 4498 123506 4510
rect 127934 4562 127986 4574
rect 127934 4498 127986 4510
rect 144174 4562 144226 4574
rect 144174 4498 144226 4510
rect 75630 4450 75682 4462
rect 22306 4398 22318 4450
rect 22370 4398 22382 4450
rect 25778 4398 25790 4450
rect 25842 4398 25854 4450
rect 28690 4398 28702 4450
rect 28754 4398 28766 4450
rect 30706 4398 30718 4450
rect 30770 4398 30782 4450
rect 34066 4398 34078 4450
rect 34130 4398 34142 4450
rect 37426 4398 37438 4450
rect 37490 4398 37502 4450
rect 41682 4398 41694 4450
rect 41746 4398 41758 4450
rect 43810 4398 43822 4450
rect 43874 4398 43886 4450
rect 45826 4398 45838 4450
rect 45890 4398 45902 4450
rect 49634 4398 49646 4450
rect 49698 4398 49710 4450
rect 52546 4398 52558 4450
rect 52610 4398 52622 4450
rect 55570 4398 55582 4450
rect 55634 4398 55646 4450
rect 57586 4398 57598 4450
rect 57650 4398 57662 4450
rect 60946 4398 60958 4450
rect 61010 4398 61022 4450
rect 67330 4398 67342 4450
rect 67394 4398 67406 4450
rect 69346 4398 69358 4450
rect 69410 4398 69422 4450
rect 73490 4398 73502 4450
rect 73554 4398 73566 4450
rect 75630 4386 75682 4398
rect 75966 4450 76018 4462
rect 75966 4386 76018 4398
rect 77422 4450 77474 4462
rect 77422 4386 77474 4398
rect 78318 4450 78370 4462
rect 78318 4386 78370 4398
rect 78878 4450 78930 4462
rect 78878 4386 78930 4398
rect 79214 4450 79266 4462
rect 79214 4386 79266 4398
rect 81678 4450 81730 4462
rect 81678 4386 81730 4398
rect 84814 4450 84866 4462
rect 84814 4386 84866 4398
rect 87838 4450 87890 4462
rect 87838 4386 87890 4398
rect 88174 4450 88226 4462
rect 88174 4386 88226 4398
rect 89294 4450 89346 4462
rect 89294 4386 89346 4398
rect 89630 4450 89682 4462
rect 89630 4386 89682 4398
rect 90190 4450 90242 4462
rect 90190 4386 90242 4398
rect 90526 4450 90578 4462
rect 90526 4386 90578 4398
rect 93998 4450 94050 4462
rect 135774 4450 135826 4462
rect 143838 4450 143890 4462
rect 94546 4398 94558 4450
rect 94610 4398 94622 4450
rect 98018 4398 98030 4450
rect 98082 4398 98094 4450
rect 101266 4398 101278 4450
rect 101330 4398 101342 4450
rect 106194 4398 106206 4450
rect 106258 4398 106270 4450
rect 107986 4398 107998 4450
rect 108050 4398 108062 4450
rect 110898 4398 110910 4450
rect 110962 4398 110974 4450
rect 113250 4398 113262 4450
rect 113314 4398 113326 4450
rect 116386 4398 116398 4450
rect 116450 4398 116462 4450
rect 119298 4398 119310 4450
rect 119362 4398 119374 4450
rect 121426 4398 121438 4450
rect 121490 4398 121502 4450
rect 124786 4398 124798 4450
rect 124850 4398 124862 4450
rect 126914 4398 126926 4450
rect 126978 4398 126990 4450
rect 129154 4398 129166 4450
rect 129218 4398 129230 4450
rect 132402 4398 132414 4450
rect 132466 4398 132478 4450
rect 134418 4398 134430 4450
rect 134482 4398 134494 4450
rect 138002 4398 138014 4450
rect 138066 4398 138078 4450
rect 140130 4398 140142 4450
rect 140194 4398 140206 4450
rect 142818 4398 142830 4450
rect 142882 4398 142894 4450
rect 146290 4398 146302 4450
rect 146354 4398 146366 4450
rect 93998 4386 94050 4398
rect 135774 4386 135826 4398
rect 143838 4386 143890 4398
rect 8878 4338 8930 4350
rect 80110 4338 80162 4350
rect 8306 4286 8318 4338
rect 8370 4286 8382 4338
rect 20066 4286 20078 4338
rect 20130 4286 20142 4338
rect 77186 4286 77198 4338
rect 77250 4286 77262 4338
rect 8878 4274 8930 4286
rect 80110 4274 80162 4286
rect 80558 4338 80610 4350
rect 104302 4338 104354 4350
rect 81442 4286 81454 4338
rect 81506 4286 81518 4338
rect 82674 4286 82686 4338
rect 82738 4286 82750 4338
rect 84578 4286 84590 4338
rect 84642 4286 84654 4338
rect 86034 4286 86046 4338
rect 86098 4286 86110 4338
rect 91074 4286 91086 4338
rect 91138 4286 91150 4338
rect 126802 4286 126814 4338
rect 126866 4286 126878 4338
rect 80558 4274 80610 4286
rect 104302 4274 104354 4286
rect 6638 4226 6690 4238
rect 15150 4226 15202 4238
rect 7186 4174 7198 4226
rect 7250 4174 7262 4226
rect 6638 4162 6690 4174
rect 15150 4162 15202 4174
rect 18286 4226 18338 4238
rect 20526 4226 20578 4238
rect 18946 4174 18958 4226
rect 19010 4174 19022 4226
rect 18286 4162 18338 4174
rect 20526 4162 20578 4174
rect 21758 4226 21810 4238
rect 25006 4226 25058 4238
rect 32958 4226 33010 4238
rect 36878 4226 36930 4238
rect 40798 4226 40850 4238
rect 48862 4226 48914 4238
rect 51998 4226 52050 4238
rect 60398 4226 60450 4238
rect 71822 4226 71874 4238
rect 23650 4174 23662 4226
rect 23714 4174 23726 4226
rect 27122 4174 27134 4226
rect 27186 4174 27198 4226
rect 30034 4174 30046 4226
rect 30098 4174 30110 4226
rect 31938 4174 31950 4226
rect 32002 4174 32014 4226
rect 35410 4174 35422 4226
rect 35474 4174 35486 4226
rect 38658 4174 38670 4226
rect 38722 4174 38734 4226
rect 43026 4174 43038 4226
rect 43090 4174 43102 4226
rect 45154 4174 45166 4226
rect 45218 4174 45230 4226
rect 47170 4174 47182 4226
rect 47234 4174 47246 4226
rect 50978 4174 50990 4226
rect 51042 4174 51054 4226
rect 53890 4174 53902 4226
rect 53954 4174 53966 4226
rect 56690 4174 56702 4226
rect 56754 4174 56766 4226
rect 58930 4174 58942 4226
rect 58994 4174 59006 4226
rect 62178 4174 62190 4226
rect 62242 4174 62254 4226
rect 68674 4174 68686 4226
rect 68738 4174 68750 4226
rect 70578 4174 70590 4226
rect 70642 4174 70654 4226
rect 21758 4162 21810 4174
rect 25006 4162 25058 4174
rect 32958 4162 33010 4174
rect 36878 4162 36930 4174
rect 40798 4162 40850 4174
rect 48862 4162 48914 4174
rect 51998 4162 52050 4174
rect 60398 4162 60450 4174
rect 71822 4162 71874 4174
rect 72606 4226 72658 4238
rect 82126 4226 82178 4238
rect 100718 4226 100770 4238
rect 103294 4226 103346 4238
rect 111806 4226 111858 4238
rect 74722 4174 74734 4226
rect 74786 4174 74798 4226
rect 83346 4174 83358 4226
rect 83410 4174 83422 4226
rect 86706 4174 86718 4226
rect 86770 4174 86782 4226
rect 91746 4174 91758 4226
rect 91810 4174 91822 4226
rect 95890 4174 95902 4226
rect 95954 4174 95966 4226
rect 99026 4174 99038 4226
rect 99090 4174 99102 4226
rect 102610 4174 102622 4226
rect 102674 4174 102686 4226
rect 103842 4174 103854 4226
rect 103906 4174 103918 4226
rect 105186 4174 105198 4226
rect 105250 4174 105262 4226
rect 109330 4174 109342 4226
rect 109394 4174 109406 4226
rect 110114 4174 110126 4226
rect 110178 4174 110190 4226
rect 72606 4162 72658 4174
rect 82126 4162 82178 4174
rect 100718 4162 100770 4174
rect 103294 4162 103346 4174
rect 111806 4162 111858 4174
rect 112254 4226 112306 4238
rect 115390 4226 115442 4238
rect 114370 4174 114382 4226
rect 114434 4174 114446 4226
rect 112254 4162 112306 4174
rect 115390 4162 115442 4174
rect 115726 4226 115778 4238
rect 124238 4226 124290 4238
rect 135326 4226 135378 4238
rect 117506 4174 117518 4226
rect 117570 4174 117582 4226
rect 118290 4174 118302 4226
rect 118354 4174 118366 4226
rect 122770 4174 122782 4226
rect 122834 4174 122846 4226
rect 125906 4174 125918 4226
rect 125970 4174 125982 4226
rect 130274 4174 130286 4226
rect 130338 4174 130350 4226
rect 131394 4174 131406 4226
rect 131458 4174 131470 4226
rect 133410 4174 133422 4226
rect 133474 4174 133486 4226
rect 115726 4162 115778 4174
rect 124238 4162 124290 4174
rect 135326 4162 135378 4174
rect 136222 4226 136274 4238
rect 139022 4226 139074 4238
rect 146862 4226 146914 4238
rect 136994 4174 137006 4226
rect 137058 4174 137070 4226
rect 141250 4174 141262 4226
rect 141314 4174 141326 4226
rect 141810 4174 141822 4226
rect 141874 4174 141886 4226
rect 144946 4174 144958 4226
rect 145010 4174 145022 4226
rect 136222 4162 136274 4174
rect 139022 4162 139074 4174
rect 146862 4162 146914 4174
rect 127598 4114 127650 4126
rect 127598 4050 127650 4062
rect 1344 3946 148624 3980
rect 1344 3894 19624 3946
rect 19676 3894 19728 3946
rect 19780 3894 19832 3946
rect 19884 3894 56444 3946
rect 56496 3894 56548 3946
rect 56600 3894 56652 3946
rect 56704 3894 93264 3946
rect 93316 3894 93368 3946
rect 93420 3894 93472 3946
rect 93524 3894 130084 3946
rect 130136 3894 130188 3946
rect 130240 3894 130292 3946
rect 130344 3894 148624 3946
rect 1344 3860 148624 3894
rect 21422 3666 21474 3678
rect 72718 3666 72770 3678
rect 86942 3666 86994 3678
rect 98590 3666 98642 3678
rect 109566 3666 109618 3678
rect 121550 3666 121602 3678
rect 126478 3666 126530 3678
rect 129278 3666 129330 3678
rect 8194 3614 8206 3666
rect 8258 3614 8270 3666
rect 10210 3614 10222 3666
rect 10274 3614 10286 3666
rect 11890 3614 11902 3666
rect 11954 3614 11966 3666
rect 19954 3614 19966 3666
rect 20018 3614 20030 3666
rect 24546 3614 24558 3666
rect 24610 3614 24622 3666
rect 28466 3614 28478 3666
rect 28530 3614 28542 3666
rect 32386 3614 32398 3666
rect 32450 3614 32462 3666
rect 36306 3614 36318 3666
rect 36370 3614 36382 3666
rect 40226 3614 40238 3666
rect 40290 3614 40302 3666
rect 43698 3614 43710 3666
rect 43762 3614 43774 3666
rect 48066 3614 48078 3666
rect 48130 3614 48142 3666
rect 51986 3614 51998 3666
rect 52050 3614 52062 3666
rect 55458 3614 55470 3666
rect 55522 3614 55534 3666
rect 59826 3614 59838 3666
rect 59890 3614 59902 3666
rect 63746 3614 63758 3666
rect 63810 3614 63822 3666
rect 67218 3614 67230 3666
rect 67282 3614 67294 3666
rect 71362 3614 71374 3666
rect 71426 3614 71438 3666
rect 75506 3614 75518 3666
rect 75570 3614 75582 3666
rect 76962 3614 76974 3666
rect 77026 3614 77038 3666
rect 78754 3614 78766 3666
rect 78818 3614 78830 3666
rect 80882 3614 80894 3666
rect 80946 3614 80958 3666
rect 82674 3614 82686 3666
rect 82738 3614 82750 3666
rect 88722 3614 88734 3666
rect 88786 3614 88798 3666
rect 90514 3614 90526 3666
rect 90578 3614 90590 3666
rect 94098 3614 94110 3666
rect 94162 3614 94174 3666
rect 97570 3614 97582 3666
rect 97634 3614 97646 3666
rect 99810 3614 99822 3666
rect 99874 3614 99886 3666
rect 103730 3614 103742 3666
rect 103794 3614 103806 3666
rect 105858 3614 105870 3666
rect 105922 3614 105934 3666
rect 107650 3614 107662 3666
rect 107714 3614 107726 3666
rect 111794 3614 111806 3666
rect 111858 3614 111870 3666
rect 116722 3614 116734 3666
rect 116786 3614 116798 3666
rect 117618 3614 117630 3666
rect 117682 3614 117694 3666
rect 119634 3614 119646 3666
rect 119698 3614 119710 3666
rect 123554 3614 123566 3666
rect 123618 3614 123630 3666
rect 128482 3614 128494 3666
rect 128546 3614 128558 3666
rect 21422 3602 21474 3614
rect 72718 3602 72770 3614
rect 86942 3602 86994 3614
rect 98590 3602 98642 3614
rect 109566 3602 109618 3614
rect 121550 3602 121602 3614
rect 126478 3602 126530 3614
rect 129278 3602 129330 3614
rect 129838 3666 129890 3678
rect 141486 3666 141538 3678
rect 131170 3614 131182 3666
rect 131234 3614 131246 3666
rect 133634 3614 133646 3666
rect 133698 3614 133710 3666
rect 135090 3614 135102 3666
rect 135154 3614 135166 3666
rect 139010 3614 139022 3666
rect 139074 3614 139086 3666
rect 143154 3614 143166 3666
rect 143218 3614 143230 3666
rect 129838 3602 129890 3614
rect 141486 3602 141538 3614
rect 30270 3554 30322 3566
rect 86494 3554 86546 3566
rect 106318 3554 106370 3566
rect 6962 3502 6974 3554
rect 7026 3502 7038 3554
rect 8754 3502 8766 3554
rect 8818 3502 8830 3554
rect 10994 3502 11006 3554
rect 11058 3502 11070 3554
rect 12786 3502 12798 3554
rect 12850 3502 12862 3554
rect 14914 3502 14926 3554
rect 14978 3502 14990 3554
rect 16706 3502 16718 3554
rect 16770 3502 16782 3554
rect 18722 3502 18734 3554
rect 18786 3502 18798 3554
rect 20626 3502 20638 3554
rect 20690 3502 20702 3554
rect 73378 3502 73390 3554
rect 73442 3502 73454 3554
rect 76290 3502 76302 3554
rect 76354 3502 76366 3554
rect 78082 3502 78094 3554
rect 78146 3502 78158 3554
rect 80210 3502 80222 3554
rect 80274 3502 80286 3554
rect 82002 3502 82014 3554
rect 82066 3502 82078 3554
rect 85362 3502 85374 3554
rect 85426 3502 85438 3554
rect 88162 3502 88174 3554
rect 88226 3502 88238 3554
rect 89842 3502 89854 3554
rect 89906 3502 89918 3554
rect 30270 3490 30322 3502
rect 86494 3490 86546 3502
rect 106318 3490 106370 3502
rect 106766 3554 106818 3566
rect 106766 3490 106818 3502
rect 110350 3554 110402 3566
rect 110350 3490 110402 3502
rect 113486 3554 113538 3566
rect 113486 3490 113538 3502
rect 118078 3554 118130 3566
rect 137006 3554 137058 3566
rect 133298 3502 133310 3554
rect 133362 3502 133374 3554
rect 118078 3490 118130 3502
rect 137006 3490 137058 3502
rect 137902 3554 137954 3566
rect 137902 3490 137954 3502
rect 25230 3442 25282 3454
rect 29150 3442 29202 3454
rect 33070 3442 33122 3454
rect 36990 3442 37042 3454
rect 40910 3442 40962 3454
rect 5842 3390 5854 3442
rect 5906 3390 5918 3442
rect 13794 3390 13806 3442
rect 13858 3390 13870 3442
rect 15586 3390 15598 3442
rect 15650 3390 15662 3442
rect 17602 3390 17614 3442
rect 17666 3390 17678 3442
rect 23426 3390 23438 3442
rect 23490 3390 23502 3442
rect 27122 3390 27134 3442
rect 27186 3390 27198 3442
rect 31378 3390 31390 3442
rect 31442 3390 31454 3442
rect 35186 3390 35198 3442
rect 35250 3390 35262 3442
rect 38882 3390 38894 3442
rect 38946 3390 38958 3442
rect 25230 3378 25282 3390
rect 29150 3378 29202 3390
rect 33070 3378 33122 3390
rect 36990 3378 37042 3390
rect 40910 3378 40962 3390
rect 41918 3442 41970 3454
rect 45390 3442 45442 3454
rect 48750 3442 48802 3454
rect 52670 3442 52722 3454
rect 42466 3390 42478 3442
rect 42530 3390 42542 3442
rect 46946 3390 46958 3442
rect 47010 3390 47022 3442
rect 50642 3390 50654 3442
rect 50706 3390 50718 3442
rect 41918 3378 41970 3390
rect 45390 3378 45442 3390
rect 48750 3378 48802 3390
rect 52670 3378 52722 3390
rect 53678 3442 53730 3454
rect 57262 3442 57314 3454
rect 60510 3442 60562 3454
rect 64430 3442 64482 3454
rect 54226 3390 54238 3442
rect 54290 3390 54302 3442
rect 58706 3390 58718 3442
rect 58770 3390 58782 3442
rect 62402 3390 62414 3442
rect 62466 3390 62478 3442
rect 53678 3378 53730 3390
rect 57262 3378 57314 3390
rect 60510 3378 60562 3390
rect 64430 3378 64482 3390
rect 65438 3442 65490 3454
rect 68910 3442 68962 3454
rect 92318 3442 92370 3454
rect 95230 3442 95282 3454
rect 98030 3442 98082 3454
rect 65986 3390 65998 3442
rect 66050 3390 66062 3442
rect 70578 3390 70590 3442
rect 70642 3390 70654 3442
rect 74498 3390 74510 3442
rect 74562 3390 74574 3442
rect 84466 3390 84478 3442
rect 84530 3390 84542 3442
rect 92866 3390 92878 3442
rect 92930 3390 92942 3442
rect 96226 3390 96238 3442
rect 96290 3390 96302 3442
rect 65438 3378 65490 3390
rect 68910 3378 68962 3390
rect 92318 3378 92370 3390
rect 95230 3378 95282 3390
rect 98030 3378 98082 3390
rect 99150 3442 99202 3454
rect 103070 3442 103122 3454
rect 113934 3442 113986 3454
rect 100818 3390 100830 3442
rect 100882 3390 100894 3442
rect 104738 3390 104750 3442
rect 104802 3390 104814 3442
rect 108658 3390 108670 3442
rect 108722 3390 108734 3442
rect 112578 3390 112590 3442
rect 112642 3390 112654 3442
rect 99150 3378 99202 3390
rect 103070 3378 103122 3390
rect 113934 3378 113986 3390
rect 114830 3442 114882 3454
rect 118526 3442 118578 3454
rect 121998 3442 122050 3454
rect 115602 3390 115614 3442
rect 115666 3390 115678 3442
rect 120642 3390 120654 3442
rect 120706 3390 120718 3442
rect 114830 3378 114882 3390
rect 118526 3378 118578 3390
rect 121998 3378 122050 3390
rect 122670 3442 122722 3454
rect 126030 3442 126082 3454
rect 130398 3442 130450 3454
rect 134206 3442 134258 3454
rect 140926 3442 140978 3454
rect 124338 3390 124350 3442
rect 124402 3390 124414 3442
rect 127362 3390 127374 3442
rect 127426 3390 127438 3442
rect 132178 3390 132190 3442
rect 132242 3390 132254 3442
rect 136098 3390 136110 3442
rect 136162 3390 136174 3442
rect 140018 3390 140030 3442
rect 140082 3390 140094 3442
rect 122670 3378 122722 3390
rect 126030 3378 126082 3390
rect 130398 3378 130450 3390
rect 134206 3378 134258 3390
rect 140926 3378 140978 3390
rect 141822 3442 141874 3454
rect 145070 3442 145122 3454
rect 144162 3390 144174 3442
rect 144226 3390 144238 3442
rect 141822 3378 141874 3390
rect 145070 3378 145122 3390
rect 73166 3330 73218 3342
rect 73166 3266 73218 3278
rect 86158 3330 86210 3342
rect 86158 3266 86210 3278
rect 110686 3330 110738 3342
rect 110686 3266 110738 3278
rect 138238 3330 138290 3342
rect 138238 3266 138290 3278
rect 1344 3162 148784 3196
rect 1344 3110 38034 3162
rect 38086 3110 38138 3162
rect 38190 3110 38242 3162
rect 38294 3110 74854 3162
rect 74906 3110 74958 3162
rect 75010 3110 75062 3162
rect 75114 3110 111674 3162
rect 111726 3110 111778 3162
rect 111830 3110 111882 3162
rect 111934 3110 148494 3162
rect 148546 3110 148598 3162
rect 148650 3110 148702 3162
rect 148754 3110 148784 3162
rect 1344 3076 148784 3110
<< via1 >>
rect 19624 36822 19676 36874
rect 19728 36822 19780 36874
rect 19832 36822 19884 36874
rect 56444 36822 56496 36874
rect 56548 36822 56600 36874
rect 56652 36822 56704 36874
rect 93264 36822 93316 36874
rect 93368 36822 93420 36874
rect 93472 36822 93524 36874
rect 130084 36822 130136 36874
rect 130188 36822 130240 36874
rect 130292 36822 130344 36874
rect 144174 36542 144226 36594
rect 147758 36542 147810 36594
rect 143054 36430 143106 36482
rect 144846 36430 144898 36482
rect 147086 36430 147138 36482
rect 145966 36318 146018 36370
rect 142158 36206 142210 36258
rect 38034 36038 38086 36090
rect 38138 36038 38190 36090
rect 38242 36038 38294 36090
rect 74854 36038 74906 36090
rect 74958 36038 75010 36090
rect 75062 36038 75114 36090
rect 111674 36038 111726 36090
rect 111778 36038 111830 36090
rect 111882 36038 111934 36090
rect 148494 36038 148546 36090
rect 148598 36038 148650 36090
rect 148702 36038 148754 36090
rect 144958 35646 145010 35698
rect 146750 35646 146802 35698
rect 143838 35534 143890 35586
rect 144286 35534 144338 35586
rect 146078 35534 146130 35586
rect 147646 35534 147698 35586
rect 19624 35254 19676 35306
rect 19728 35254 19780 35306
rect 19832 35254 19884 35306
rect 56444 35254 56496 35306
rect 56548 35254 56600 35306
rect 56652 35254 56704 35306
rect 93264 35254 93316 35306
rect 93368 35254 93420 35306
rect 93472 35254 93524 35306
rect 130084 35254 130136 35306
rect 130188 35254 130240 35306
rect 130292 35254 130344 35306
rect 144958 34862 145010 34914
rect 146078 34750 146130 34802
rect 144398 34638 144450 34690
rect 146638 34638 146690 34690
rect 147086 34638 147138 34690
rect 38034 34470 38086 34522
rect 38138 34470 38190 34522
rect 38242 34470 38294 34522
rect 74854 34470 74906 34522
rect 74958 34470 75010 34522
rect 75062 34470 75114 34522
rect 111674 34470 111726 34522
rect 111778 34470 111830 34522
rect 111882 34470 111934 34522
rect 148494 34470 148546 34522
rect 148598 34470 148650 34522
rect 148702 34470 148754 34522
rect 144958 34078 145010 34130
rect 144286 33966 144338 34018
rect 146078 33966 146130 34018
rect 19624 33686 19676 33738
rect 19728 33686 19780 33738
rect 19832 33686 19884 33738
rect 56444 33686 56496 33738
rect 56548 33686 56600 33738
rect 56652 33686 56704 33738
rect 93264 33686 93316 33738
rect 93368 33686 93420 33738
rect 93472 33686 93524 33738
rect 130084 33686 130136 33738
rect 130188 33686 130240 33738
rect 130292 33686 130344 33738
rect 144958 33294 145010 33346
rect 146078 33182 146130 33234
rect 144398 33070 144450 33122
rect 38034 32902 38086 32954
rect 38138 32902 38190 32954
rect 38242 32902 38294 32954
rect 74854 32902 74906 32954
rect 74958 32902 75010 32954
rect 75062 32902 75114 32954
rect 111674 32902 111726 32954
rect 111778 32902 111830 32954
rect 111882 32902 111934 32954
rect 148494 32902 148546 32954
rect 148598 32902 148650 32954
rect 148702 32902 148754 32954
rect 19624 32118 19676 32170
rect 19728 32118 19780 32170
rect 19832 32118 19884 32170
rect 56444 32118 56496 32170
rect 56548 32118 56600 32170
rect 56652 32118 56704 32170
rect 93264 32118 93316 32170
rect 93368 32118 93420 32170
rect 93472 32118 93524 32170
rect 130084 32118 130136 32170
rect 130188 32118 130240 32170
rect 130292 32118 130344 32170
rect 144958 31726 145010 31778
rect 146078 31614 146130 31666
rect 144398 31502 144450 31554
rect 38034 31334 38086 31386
rect 38138 31334 38190 31386
rect 38242 31334 38294 31386
rect 74854 31334 74906 31386
rect 74958 31334 75010 31386
rect 75062 31334 75114 31386
rect 111674 31334 111726 31386
rect 111778 31334 111830 31386
rect 111882 31334 111934 31386
rect 148494 31334 148546 31386
rect 148598 31334 148650 31386
rect 148702 31334 148754 31386
rect 144958 30942 145010 30994
rect 144286 30830 144338 30882
rect 146078 30830 146130 30882
rect 19624 30550 19676 30602
rect 19728 30550 19780 30602
rect 19832 30550 19884 30602
rect 56444 30550 56496 30602
rect 56548 30550 56600 30602
rect 56652 30550 56704 30602
rect 93264 30550 93316 30602
rect 93368 30550 93420 30602
rect 93472 30550 93524 30602
rect 130084 30550 130136 30602
rect 130188 30550 130240 30602
rect 130292 30550 130344 30602
rect 144958 30158 145010 30210
rect 146078 30046 146130 30098
rect 144398 29934 144450 29986
rect 38034 29766 38086 29818
rect 38138 29766 38190 29818
rect 38242 29766 38294 29818
rect 74854 29766 74906 29818
rect 74958 29766 75010 29818
rect 75062 29766 75114 29818
rect 111674 29766 111726 29818
rect 111778 29766 111830 29818
rect 111882 29766 111934 29818
rect 148494 29766 148546 29818
rect 148598 29766 148650 29818
rect 148702 29766 148754 29818
rect 144958 29374 145010 29426
rect 144286 29262 144338 29314
rect 146078 29262 146130 29314
rect 19624 28982 19676 29034
rect 19728 28982 19780 29034
rect 19832 28982 19884 29034
rect 56444 28982 56496 29034
rect 56548 28982 56600 29034
rect 56652 28982 56704 29034
rect 93264 28982 93316 29034
rect 93368 28982 93420 29034
rect 93472 28982 93524 29034
rect 130084 28982 130136 29034
rect 130188 28982 130240 29034
rect 130292 28982 130344 29034
rect 144398 28590 144450 28642
rect 144958 28590 145010 28642
rect 146078 28590 146130 28642
rect 38034 28198 38086 28250
rect 38138 28198 38190 28250
rect 38242 28198 38294 28250
rect 74854 28198 74906 28250
rect 74958 28198 75010 28250
rect 75062 28198 75114 28250
rect 111674 28198 111726 28250
rect 111778 28198 111830 28250
rect 111882 28198 111934 28250
rect 148494 28198 148546 28250
rect 148598 28198 148650 28250
rect 148702 28198 148754 28250
rect 144958 27806 145010 27858
rect 144286 27694 144338 27746
rect 146078 27694 146130 27746
rect 19624 27414 19676 27466
rect 19728 27414 19780 27466
rect 19832 27414 19884 27466
rect 56444 27414 56496 27466
rect 56548 27414 56600 27466
rect 56652 27414 56704 27466
rect 93264 27414 93316 27466
rect 93368 27414 93420 27466
rect 93472 27414 93524 27466
rect 130084 27414 130136 27466
rect 130188 27414 130240 27466
rect 130292 27414 130344 27466
rect 144958 27022 145010 27074
rect 144398 26910 144450 26962
rect 146078 26910 146130 26962
rect 38034 26630 38086 26682
rect 38138 26630 38190 26682
rect 38242 26630 38294 26682
rect 74854 26630 74906 26682
rect 74958 26630 75010 26682
rect 75062 26630 75114 26682
rect 111674 26630 111726 26682
rect 111778 26630 111830 26682
rect 111882 26630 111934 26682
rect 148494 26630 148546 26682
rect 148598 26630 148650 26682
rect 148702 26630 148754 26682
rect 19624 25846 19676 25898
rect 19728 25846 19780 25898
rect 19832 25846 19884 25898
rect 56444 25846 56496 25898
rect 56548 25846 56600 25898
rect 56652 25846 56704 25898
rect 93264 25846 93316 25898
rect 93368 25846 93420 25898
rect 93472 25846 93524 25898
rect 130084 25846 130136 25898
rect 130188 25846 130240 25898
rect 130292 25846 130344 25898
rect 144958 25454 145010 25506
rect 146078 25342 146130 25394
rect 144398 25230 144450 25282
rect 38034 25062 38086 25114
rect 38138 25062 38190 25114
rect 38242 25062 38294 25114
rect 74854 25062 74906 25114
rect 74958 25062 75010 25114
rect 75062 25062 75114 25114
rect 111674 25062 111726 25114
rect 111778 25062 111830 25114
rect 111882 25062 111934 25114
rect 148494 25062 148546 25114
rect 148598 25062 148650 25114
rect 148702 25062 148754 25114
rect 144958 24670 145010 24722
rect 144286 24558 144338 24610
rect 146078 24558 146130 24610
rect 19624 24278 19676 24330
rect 19728 24278 19780 24330
rect 19832 24278 19884 24330
rect 56444 24278 56496 24330
rect 56548 24278 56600 24330
rect 56652 24278 56704 24330
rect 93264 24278 93316 24330
rect 93368 24278 93420 24330
rect 93472 24278 93524 24330
rect 130084 24278 130136 24330
rect 130188 24278 130240 24330
rect 130292 24278 130344 24330
rect 144958 23886 145010 23938
rect 146078 23774 146130 23826
rect 144398 23662 144450 23714
rect 38034 23494 38086 23546
rect 38138 23494 38190 23546
rect 38242 23494 38294 23546
rect 74854 23494 74906 23546
rect 74958 23494 75010 23546
rect 75062 23494 75114 23546
rect 111674 23494 111726 23546
rect 111778 23494 111830 23546
rect 111882 23494 111934 23546
rect 148494 23494 148546 23546
rect 148598 23494 148650 23546
rect 148702 23494 148754 23546
rect 144958 23102 145010 23154
rect 144286 22990 144338 23042
rect 146078 22990 146130 23042
rect 19624 22710 19676 22762
rect 19728 22710 19780 22762
rect 19832 22710 19884 22762
rect 56444 22710 56496 22762
rect 56548 22710 56600 22762
rect 56652 22710 56704 22762
rect 93264 22710 93316 22762
rect 93368 22710 93420 22762
rect 93472 22710 93524 22762
rect 130084 22710 130136 22762
rect 130188 22710 130240 22762
rect 130292 22710 130344 22762
rect 144958 22318 145010 22370
rect 146078 22206 146130 22258
rect 144398 22094 144450 22146
rect 38034 21926 38086 21978
rect 38138 21926 38190 21978
rect 38242 21926 38294 21978
rect 74854 21926 74906 21978
rect 74958 21926 75010 21978
rect 75062 21926 75114 21978
rect 111674 21926 111726 21978
rect 111778 21926 111830 21978
rect 111882 21926 111934 21978
rect 148494 21926 148546 21978
rect 148598 21926 148650 21978
rect 148702 21926 148754 21978
rect 144958 21534 145010 21586
rect 144286 21422 144338 21474
rect 146078 21422 146130 21474
rect 19624 21142 19676 21194
rect 19728 21142 19780 21194
rect 19832 21142 19884 21194
rect 56444 21142 56496 21194
rect 56548 21142 56600 21194
rect 56652 21142 56704 21194
rect 93264 21142 93316 21194
rect 93368 21142 93420 21194
rect 93472 21142 93524 21194
rect 130084 21142 130136 21194
rect 130188 21142 130240 21194
rect 130292 21142 130344 21194
rect 144958 20750 145010 20802
rect 146078 20638 146130 20690
rect 144398 20526 144450 20578
rect 38034 20358 38086 20410
rect 38138 20358 38190 20410
rect 38242 20358 38294 20410
rect 74854 20358 74906 20410
rect 74958 20358 75010 20410
rect 75062 20358 75114 20410
rect 111674 20358 111726 20410
rect 111778 20358 111830 20410
rect 111882 20358 111934 20410
rect 148494 20358 148546 20410
rect 148598 20358 148650 20410
rect 148702 20358 148754 20410
rect 19624 19574 19676 19626
rect 19728 19574 19780 19626
rect 19832 19574 19884 19626
rect 56444 19574 56496 19626
rect 56548 19574 56600 19626
rect 56652 19574 56704 19626
rect 93264 19574 93316 19626
rect 93368 19574 93420 19626
rect 93472 19574 93524 19626
rect 130084 19574 130136 19626
rect 130188 19574 130240 19626
rect 130292 19574 130344 19626
rect 144958 19182 145010 19234
rect 146078 19070 146130 19122
rect 144398 18958 144450 19010
rect 38034 18790 38086 18842
rect 38138 18790 38190 18842
rect 38242 18790 38294 18842
rect 74854 18790 74906 18842
rect 74958 18790 75010 18842
rect 75062 18790 75114 18842
rect 111674 18790 111726 18842
rect 111778 18790 111830 18842
rect 111882 18790 111934 18842
rect 148494 18790 148546 18842
rect 148598 18790 148650 18842
rect 148702 18790 148754 18842
rect 111582 18622 111634 18674
rect 111246 18510 111298 18562
rect 144958 18398 145010 18450
rect 110686 18286 110738 18338
rect 144286 18286 144338 18338
rect 146078 18286 146130 18338
rect 19624 18006 19676 18058
rect 19728 18006 19780 18058
rect 19832 18006 19884 18058
rect 56444 18006 56496 18058
rect 56548 18006 56600 18058
rect 56652 18006 56704 18058
rect 93264 18006 93316 18058
rect 93368 18006 93420 18058
rect 93472 18006 93524 18058
rect 130084 18006 130136 18058
rect 130188 18006 130240 18058
rect 130292 18006 130344 18058
rect 144958 17614 145010 17666
rect 146078 17502 146130 17554
rect 144398 17390 144450 17442
rect 38034 17222 38086 17274
rect 38138 17222 38190 17274
rect 38242 17222 38294 17274
rect 74854 17222 74906 17274
rect 74958 17222 75010 17274
rect 75062 17222 75114 17274
rect 111674 17222 111726 17274
rect 111778 17222 111830 17274
rect 111882 17222 111934 17274
rect 148494 17222 148546 17274
rect 148598 17222 148650 17274
rect 148702 17222 148754 17274
rect 144286 16830 144338 16882
rect 144958 16830 145010 16882
rect 146078 16830 146130 16882
rect 19624 16438 19676 16490
rect 19728 16438 19780 16490
rect 19832 16438 19884 16490
rect 56444 16438 56496 16490
rect 56548 16438 56600 16490
rect 56652 16438 56704 16490
rect 93264 16438 93316 16490
rect 93368 16438 93420 16490
rect 93472 16438 93524 16490
rect 130084 16438 130136 16490
rect 130188 16438 130240 16490
rect 130292 16438 130344 16490
rect 144958 16046 145010 16098
rect 146078 15934 146130 15986
rect 144398 15822 144450 15874
rect 38034 15654 38086 15706
rect 38138 15654 38190 15706
rect 38242 15654 38294 15706
rect 74854 15654 74906 15706
rect 74958 15654 75010 15706
rect 75062 15654 75114 15706
rect 111674 15654 111726 15706
rect 111778 15654 111830 15706
rect 111882 15654 111934 15706
rect 148494 15654 148546 15706
rect 148598 15654 148650 15706
rect 148702 15654 148754 15706
rect 144958 15262 145010 15314
rect 144286 15150 144338 15202
rect 146078 15150 146130 15202
rect 19624 14870 19676 14922
rect 19728 14870 19780 14922
rect 19832 14870 19884 14922
rect 56444 14870 56496 14922
rect 56548 14870 56600 14922
rect 56652 14870 56704 14922
rect 93264 14870 93316 14922
rect 93368 14870 93420 14922
rect 93472 14870 93524 14922
rect 130084 14870 130136 14922
rect 130188 14870 130240 14922
rect 130292 14870 130344 14922
rect 144958 14478 145010 14530
rect 146078 14366 146130 14418
rect 144398 14254 144450 14306
rect 38034 14086 38086 14138
rect 38138 14086 38190 14138
rect 38242 14086 38294 14138
rect 74854 14086 74906 14138
rect 74958 14086 75010 14138
rect 75062 14086 75114 14138
rect 111674 14086 111726 14138
rect 111778 14086 111830 14138
rect 111882 14086 111934 14138
rect 148494 14086 148546 14138
rect 148598 14086 148650 14138
rect 148702 14086 148754 14138
rect 19624 13302 19676 13354
rect 19728 13302 19780 13354
rect 19832 13302 19884 13354
rect 56444 13302 56496 13354
rect 56548 13302 56600 13354
rect 56652 13302 56704 13354
rect 93264 13302 93316 13354
rect 93368 13302 93420 13354
rect 93472 13302 93524 13354
rect 130084 13302 130136 13354
rect 130188 13302 130240 13354
rect 130292 13302 130344 13354
rect 144958 12910 145010 12962
rect 101166 12798 101218 12850
rect 101502 12798 101554 12850
rect 146078 12798 146130 12850
rect 144398 12686 144450 12738
rect 38034 12518 38086 12570
rect 38138 12518 38190 12570
rect 38242 12518 38294 12570
rect 74854 12518 74906 12570
rect 74958 12518 75010 12570
rect 75062 12518 75114 12570
rect 111674 12518 111726 12570
rect 111778 12518 111830 12570
rect 111882 12518 111934 12570
rect 148494 12518 148546 12570
rect 148598 12518 148650 12570
rect 148702 12518 148754 12570
rect 100494 12350 100546 12402
rect 100158 12126 100210 12178
rect 144958 12126 145010 12178
rect 144286 12014 144338 12066
rect 146078 12014 146130 12066
rect 19624 11734 19676 11786
rect 19728 11734 19780 11786
rect 19832 11734 19884 11786
rect 56444 11734 56496 11786
rect 56548 11734 56600 11786
rect 56652 11734 56704 11786
rect 93264 11734 93316 11786
rect 93368 11734 93420 11786
rect 93472 11734 93524 11786
rect 130084 11734 130136 11786
rect 130188 11734 130240 11786
rect 130292 11734 130344 11786
rect 144958 11342 145010 11394
rect 101166 11230 101218 11282
rect 146078 11230 146130 11282
rect 100494 11118 100546 11170
rect 101502 11118 101554 11170
rect 144398 11118 144450 11170
rect 38034 10950 38086 11002
rect 38138 10950 38190 11002
rect 38242 10950 38294 11002
rect 74854 10950 74906 11002
rect 74958 10950 75010 11002
rect 75062 10950 75114 11002
rect 111674 10950 111726 11002
rect 111778 10950 111830 11002
rect 111882 10950 111934 11002
rect 148494 10950 148546 11002
rect 148598 10950 148650 11002
rect 148702 10950 148754 11002
rect 146302 10670 146354 10722
rect 145182 10446 145234 10498
rect 146862 10446 146914 10498
rect 19624 10166 19676 10218
rect 19728 10166 19780 10218
rect 19832 10166 19884 10218
rect 56444 10166 56496 10218
rect 56548 10166 56600 10218
rect 56652 10166 56704 10218
rect 93264 10166 93316 10218
rect 93368 10166 93420 10218
rect 93472 10166 93524 10218
rect 130084 10166 130136 10218
rect 130188 10166 130240 10218
rect 130292 10166 130344 10218
rect 144958 9886 145010 9938
rect 146302 9662 146354 9714
rect 146974 9550 147026 9602
rect 38034 9382 38086 9434
rect 38138 9382 38190 9434
rect 38242 9382 38294 9434
rect 74854 9382 74906 9434
rect 74958 9382 75010 9434
rect 75062 9382 75114 9434
rect 111674 9382 111726 9434
rect 111778 9382 111830 9434
rect 111882 9382 111934 9434
rect 148494 9382 148546 9434
rect 148598 9382 148650 9434
rect 148702 9382 148754 9434
rect 146302 9102 146354 9154
rect 144958 8878 145010 8930
rect 146862 8878 146914 8930
rect 19624 8598 19676 8650
rect 19728 8598 19780 8650
rect 19832 8598 19884 8650
rect 56444 8598 56496 8650
rect 56548 8598 56600 8650
rect 56652 8598 56704 8650
rect 93264 8598 93316 8650
rect 93368 8598 93420 8650
rect 93472 8598 93524 8650
rect 130084 8598 130136 8650
rect 130188 8598 130240 8650
rect 130292 8598 130344 8650
rect 144958 8318 145010 8370
rect 146302 8094 146354 8146
rect 146974 7982 147026 8034
rect 38034 7814 38086 7866
rect 38138 7814 38190 7866
rect 38242 7814 38294 7866
rect 74854 7814 74906 7866
rect 74958 7814 75010 7866
rect 75062 7814 75114 7866
rect 111674 7814 111726 7866
rect 111778 7814 111830 7866
rect 111882 7814 111934 7866
rect 148494 7814 148546 7866
rect 148598 7814 148650 7866
rect 148702 7814 148754 7866
rect 105534 7646 105586 7698
rect 139022 7646 139074 7698
rect 139918 7646 139970 7698
rect 129838 7534 129890 7586
rect 130958 7534 131010 7586
rect 131294 7534 131346 7586
rect 131742 7534 131794 7586
rect 146190 7534 146242 7586
rect 146862 7534 146914 7586
rect 105310 7422 105362 7474
rect 138798 7422 138850 7474
rect 139694 7422 139746 7474
rect 130398 7310 130450 7362
rect 137790 7310 137842 7362
rect 140366 7310 140418 7362
rect 144286 7310 144338 7362
rect 144958 7310 145010 7362
rect 130398 7198 130450 7250
rect 130622 7198 130674 7250
rect 19624 7030 19676 7082
rect 19728 7030 19780 7082
rect 19832 7030 19884 7082
rect 56444 7030 56496 7082
rect 56548 7030 56600 7082
rect 56652 7030 56704 7082
rect 93264 7030 93316 7082
rect 93368 7030 93420 7082
rect 93472 7030 93524 7082
rect 130084 7030 130136 7082
rect 130188 7030 130240 7082
rect 130292 7030 130344 7082
rect 139246 6862 139298 6914
rect 138910 6750 138962 6802
rect 142942 6750 142994 6802
rect 145070 6750 145122 6802
rect 110462 6638 110514 6690
rect 117966 6638 118018 6690
rect 128830 6638 128882 6690
rect 129614 6638 129666 6690
rect 131966 6638 132018 6690
rect 137566 6638 137618 6690
rect 139918 6638 139970 6690
rect 101166 6526 101218 6578
rect 101502 6526 101554 6578
rect 103294 6526 103346 6578
rect 103630 6526 103682 6578
rect 104190 6526 104242 6578
rect 104526 6526 104578 6578
rect 105198 6526 105250 6578
rect 105534 6526 105586 6578
rect 117070 6526 117122 6578
rect 117406 6526 117458 6578
rect 130174 6526 130226 6578
rect 130510 6526 130562 6578
rect 131070 6526 131122 6578
rect 131406 6526 131458 6578
rect 132974 6526 133026 6578
rect 133310 6526 133362 6578
rect 138126 6526 138178 6578
rect 138686 6526 138738 6578
rect 140926 6526 140978 6578
rect 141262 6526 141314 6578
rect 144286 6526 144338 6578
rect 146302 6526 146354 6578
rect 146974 6526 147026 6578
rect 105982 6414 106034 6466
rect 111022 6414 111074 6466
rect 111470 6414 111522 6466
rect 112702 6414 112754 6466
rect 124350 6414 124402 6466
rect 129278 6414 129330 6466
rect 133982 6414 134034 6466
rect 137006 6414 137058 6466
rect 38034 6246 38086 6298
rect 38138 6246 38190 6298
rect 38242 6246 38294 6298
rect 74854 6246 74906 6298
rect 74958 6246 75010 6298
rect 75062 6246 75114 6298
rect 111674 6246 111726 6298
rect 111778 6246 111830 6298
rect 111882 6246 111934 6298
rect 148494 6246 148546 6298
rect 148598 6246 148650 6298
rect 148702 6246 148754 6298
rect 82798 6078 82850 6130
rect 86942 6078 86994 6130
rect 88398 6078 88450 6130
rect 98478 6078 98530 6130
rect 101950 6078 102002 6130
rect 103742 6078 103794 6130
rect 105310 6078 105362 6130
rect 106990 6078 107042 6130
rect 109118 6078 109170 6130
rect 110910 6078 110962 6130
rect 113486 6078 113538 6130
rect 115278 6078 115330 6130
rect 120094 6078 120146 6130
rect 122110 6078 122162 6130
rect 124910 6078 124962 6130
rect 126030 6078 126082 6130
rect 130510 6078 130562 6130
rect 134766 6078 134818 6130
rect 136222 6078 136274 6130
rect 137342 6078 137394 6130
rect 141150 6078 141202 6130
rect 142158 6078 142210 6130
rect 97470 5966 97522 6018
rect 97918 5966 97970 6018
rect 102734 5966 102786 6018
rect 106206 5966 106258 6018
rect 109902 5966 109954 6018
rect 112030 5966 112082 6018
rect 116062 5966 116114 6018
rect 116510 5966 116562 6018
rect 118078 5966 118130 6018
rect 122894 5966 122946 6018
rect 123342 5966 123394 6018
rect 129502 5966 129554 6018
rect 129950 5966 130002 6018
rect 131742 5966 131794 6018
rect 132078 5966 132130 6018
rect 138238 5966 138290 6018
rect 138686 5966 138738 6018
rect 140142 5966 140194 6018
rect 144062 5966 144114 6018
rect 146302 5966 146354 6018
rect 102622 5854 102674 5906
rect 106430 5854 106482 5906
rect 109790 5854 109842 5906
rect 111806 5854 111858 5906
rect 113262 5854 113314 5906
rect 117966 5854 118018 5906
rect 119086 5854 119138 5906
rect 119758 5854 119810 5906
rect 123902 5854 123954 5906
rect 124574 5854 124626 5906
rect 125806 5854 125858 5906
rect 132638 5854 132690 5906
rect 133310 5854 133362 5906
rect 134430 5854 134482 5906
rect 137006 5854 137058 5906
rect 140366 5854 140418 5906
rect 141822 5854 141874 5906
rect 75742 5742 75794 5794
rect 86046 5742 86098 5794
rect 96462 5742 96514 5794
rect 99038 5742 99090 5794
rect 99486 5742 99538 5794
rect 101502 5742 101554 5794
rect 104414 5742 104466 5794
rect 107438 5742 107490 5794
rect 107886 5742 107938 5794
rect 108782 5742 108834 5794
rect 114718 5742 114770 5794
rect 126590 5742 126642 5794
rect 127822 5742 127874 5794
rect 128270 5742 128322 5794
rect 133758 5742 133810 5794
rect 135886 5742 135938 5794
rect 142718 5742 142770 5794
rect 144958 5742 145010 5794
rect 146862 5742 146914 5794
rect 147310 5742 147362 5794
rect 98142 5630 98194 5682
rect 103406 5630 103458 5682
rect 105646 5630 105698 5682
rect 106766 5630 106818 5682
rect 107438 5630 107490 5682
rect 110574 5630 110626 5682
rect 116734 5630 116786 5682
rect 117070 5630 117122 5682
rect 118750 5630 118802 5682
rect 123566 5630 123618 5682
rect 130174 5630 130226 5682
rect 132302 5630 132354 5682
rect 138910 5630 138962 5682
rect 139246 5630 139298 5682
rect 140814 5630 140866 5682
rect 19624 5462 19676 5514
rect 19728 5462 19780 5514
rect 19832 5462 19884 5514
rect 56444 5462 56496 5514
rect 56548 5462 56600 5514
rect 56652 5462 56704 5514
rect 93264 5462 93316 5514
rect 93368 5462 93420 5514
rect 93472 5462 93524 5514
rect 130084 5462 130136 5514
rect 130188 5462 130240 5514
rect 130292 5462 130344 5514
rect 96238 5294 96290 5346
rect 98142 5294 98194 5346
rect 100046 5294 100098 5346
rect 102958 5294 103010 5346
rect 104862 5294 104914 5346
rect 112254 5294 112306 5346
rect 114158 5294 114210 5346
rect 116174 5294 116226 5346
rect 126254 5294 126306 5346
rect 129726 5294 129778 5346
rect 131742 5294 131794 5346
rect 135438 5294 135490 5346
rect 137342 5294 137394 5346
rect 139246 5294 139298 5346
rect 65662 5182 65714 5234
rect 76190 5182 76242 5234
rect 77646 5182 77698 5234
rect 79438 5182 79490 5234
rect 89854 5182 89906 5234
rect 90302 5182 90354 5234
rect 90750 5182 90802 5234
rect 142942 5182 142994 5234
rect 144958 5182 145010 5234
rect 63758 5070 63810 5122
rect 78542 5070 78594 5122
rect 81006 5070 81058 5122
rect 81454 5070 81506 5122
rect 82238 5070 82290 5122
rect 83358 5070 83410 5122
rect 83806 5070 83858 5122
rect 86718 5070 86770 5122
rect 89406 5070 89458 5122
rect 95454 5070 95506 5122
rect 95902 5070 95954 5122
rect 97358 5070 97410 5122
rect 97806 5070 97858 5122
rect 99262 5070 99314 5122
rect 99710 5070 99762 5122
rect 101054 5070 101106 5122
rect 102174 5070 102226 5122
rect 102622 5070 102674 5122
rect 103742 5070 103794 5122
rect 104526 5070 104578 5122
rect 105870 5070 105922 5122
rect 106430 5070 106482 5122
rect 109566 5070 109618 5122
rect 110014 5070 110066 5122
rect 111470 5070 111522 5122
rect 111918 5070 111970 5122
rect 113150 5070 113202 5122
rect 113822 5070 113874 5122
rect 115390 5070 115442 5122
rect 115838 5070 115890 5122
rect 117966 5070 118018 5122
rect 122334 5070 122386 5122
rect 122782 5070 122834 5122
rect 125470 5070 125522 5122
rect 125918 5070 125970 5122
rect 128942 5070 128994 5122
rect 129390 5070 129442 5122
rect 130958 5070 131010 5122
rect 131406 5070 131458 5122
rect 133534 5070 133586 5122
rect 134654 5070 134706 5122
rect 135102 5070 135154 5122
rect 136558 5070 136610 5122
rect 137006 5070 137058 5122
rect 138462 5070 138514 5122
rect 138910 5070 138962 5122
rect 139806 5070 139858 5122
rect 141150 5070 141202 5122
rect 141822 5070 141874 5122
rect 146862 5070 146914 5122
rect 64318 4958 64370 5010
rect 75406 4958 75458 5010
rect 80670 4958 80722 5010
rect 85486 4958 85538 5010
rect 87726 4958 87778 5010
rect 95118 4958 95170 5010
rect 97022 4958 97074 5010
rect 98926 4958 98978 5010
rect 101838 4958 101890 5010
rect 103966 4958 104018 5010
rect 105646 4958 105698 5010
rect 106766 4958 106818 5010
rect 107438 4958 107490 5010
rect 107774 4958 107826 5010
rect 109230 4958 109282 5010
rect 111134 4958 111186 5010
rect 113038 4958 113090 5010
rect 115054 4958 115106 5010
rect 117182 4958 117234 5010
rect 117742 4958 117794 5010
rect 118302 4958 118354 5010
rect 118974 4958 119026 5010
rect 119310 4958 119362 5010
rect 119870 4958 119922 5010
rect 120206 4958 120258 5010
rect 121998 4958 122050 5010
rect 123118 4958 123170 5010
rect 123790 4958 123842 5010
rect 124126 4958 124178 5010
rect 125134 4958 125186 5010
rect 126814 4958 126866 5010
rect 127598 4958 127650 5010
rect 127934 4958 127986 5010
rect 128830 4958 128882 5010
rect 130622 4958 130674 5010
rect 132974 4958 133026 5010
rect 134430 4958 134482 5010
rect 136446 4958 136498 5010
rect 138350 4958 138402 5010
rect 141262 4958 141314 5010
rect 144286 4958 144338 5010
rect 146302 4958 146354 5010
rect 30382 4846 30434 4898
rect 45502 4846 45554 4898
rect 56926 4846 56978 4898
rect 69358 4846 69410 4898
rect 75742 4846 75794 4898
rect 82462 4846 82514 4898
rect 83022 4846 83074 4898
rect 85822 4846 85874 4898
rect 86382 4846 86434 4898
rect 87390 4846 87442 4898
rect 88174 4846 88226 4898
rect 89070 4846 89122 4898
rect 94558 4846 94610 4898
rect 108222 4846 108274 4898
rect 110350 4846 110402 4898
rect 121438 4846 121490 4898
rect 142158 4846 142210 4898
rect 147422 4846 147474 4898
rect 38034 4678 38086 4730
rect 38138 4678 38190 4730
rect 38242 4678 38294 4730
rect 74854 4678 74906 4730
rect 74958 4678 75010 4730
rect 75062 4678 75114 4730
rect 111674 4678 111726 4730
rect 111778 4678 111830 4730
rect 111882 4678 111934 4730
rect 148494 4678 148546 4730
rect 148598 4678 148650 4730
rect 148702 4678 148754 4730
rect 9774 4510 9826 4562
rect 11342 4510 11394 4562
rect 13022 4510 13074 4562
rect 17054 4510 17106 4562
rect 76526 4510 76578 4562
rect 77982 4510 78034 4562
rect 79774 4510 79826 4562
rect 85374 4510 85426 4562
rect 96462 4510 96514 4562
rect 97134 4510 97186 4562
rect 107102 4510 107154 4562
rect 120206 4510 120258 4562
rect 123454 4510 123506 4562
rect 127934 4510 127986 4562
rect 144174 4510 144226 4562
rect 22318 4398 22370 4450
rect 25790 4398 25842 4450
rect 28702 4398 28754 4450
rect 30718 4398 30770 4450
rect 34078 4398 34130 4450
rect 37438 4398 37490 4450
rect 41694 4398 41746 4450
rect 43822 4398 43874 4450
rect 45838 4398 45890 4450
rect 49646 4398 49698 4450
rect 52558 4398 52610 4450
rect 55582 4398 55634 4450
rect 57598 4398 57650 4450
rect 60958 4398 61010 4450
rect 67342 4398 67394 4450
rect 69358 4398 69410 4450
rect 73502 4398 73554 4450
rect 75630 4398 75682 4450
rect 75966 4398 76018 4450
rect 77422 4398 77474 4450
rect 78318 4398 78370 4450
rect 78878 4398 78930 4450
rect 79214 4398 79266 4450
rect 81678 4398 81730 4450
rect 84814 4398 84866 4450
rect 87838 4398 87890 4450
rect 88174 4398 88226 4450
rect 89294 4398 89346 4450
rect 89630 4398 89682 4450
rect 90190 4398 90242 4450
rect 90526 4398 90578 4450
rect 93998 4398 94050 4450
rect 94558 4398 94610 4450
rect 98030 4398 98082 4450
rect 101278 4398 101330 4450
rect 106206 4398 106258 4450
rect 107998 4398 108050 4450
rect 110910 4398 110962 4450
rect 113262 4398 113314 4450
rect 116398 4398 116450 4450
rect 119310 4398 119362 4450
rect 121438 4398 121490 4450
rect 124798 4398 124850 4450
rect 126926 4398 126978 4450
rect 129166 4398 129218 4450
rect 132414 4398 132466 4450
rect 134430 4398 134482 4450
rect 135774 4398 135826 4450
rect 138014 4398 138066 4450
rect 140142 4398 140194 4450
rect 142830 4398 142882 4450
rect 143838 4398 143890 4450
rect 146302 4398 146354 4450
rect 8318 4286 8370 4338
rect 8878 4286 8930 4338
rect 20078 4286 20130 4338
rect 77198 4286 77250 4338
rect 80110 4286 80162 4338
rect 80558 4286 80610 4338
rect 81454 4286 81506 4338
rect 82686 4286 82738 4338
rect 84590 4286 84642 4338
rect 86046 4286 86098 4338
rect 91086 4286 91138 4338
rect 104302 4286 104354 4338
rect 126814 4286 126866 4338
rect 6638 4174 6690 4226
rect 7198 4174 7250 4226
rect 15150 4174 15202 4226
rect 18286 4174 18338 4226
rect 18958 4174 19010 4226
rect 20526 4174 20578 4226
rect 21758 4174 21810 4226
rect 23662 4174 23714 4226
rect 25006 4174 25058 4226
rect 27134 4174 27186 4226
rect 30046 4174 30098 4226
rect 31950 4174 32002 4226
rect 32958 4174 33010 4226
rect 35422 4174 35474 4226
rect 36878 4174 36930 4226
rect 38670 4174 38722 4226
rect 40798 4174 40850 4226
rect 43038 4174 43090 4226
rect 45166 4174 45218 4226
rect 47182 4174 47234 4226
rect 48862 4174 48914 4226
rect 50990 4174 51042 4226
rect 51998 4174 52050 4226
rect 53902 4174 53954 4226
rect 56702 4174 56754 4226
rect 58942 4174 58994 4226
rect 60398 4174 60450 4226
rect 62190 4174 62242 4226
rect 68686 4174 68738 4226
rect 70590 4174 70642 4226
rect 71822 4174 71874 4226
rect 72606 4174 72658 4226
rect 74734 4174 74786 4226
rect 82126 4174 82178 4226
rect 83358 4174 83410 4226
rect 86718 4174 86770 4226
rect 91758 4174 91810 4226
rect 95902 4174 95954 4226
rect 99038 4174 99090 4226
rect 100718 4174 100770 4226
rect 102622 4174 102674 4226
rect 103294 4174 103346 4226
rect 103854 4174 103906 4226
rect 105198 4174 105250 4226
rect 109342 4174 109394 4226
rect 110126 4174 110178 4226
rect 111806 4174 111858 4226
rect 112254 4174 112306 4226
rect 114382 4174 114434 4226
rect 115390 4174 115442 4226
rect 115726 4174 115778 4226
rect 117518 4174 117570 4226
rect 118302 4174 118354 4226
rect 122782 4174 122834 4226
rect 124238 4174 124290 4226
rect 125918 4174 125970 4226
rect 130286 4174 130338 4226
rect 131406 4174 131458 4226
rect 133422 4174 133474 4226
rect 135326 4174 135378 4226
rect 136222 4174 136274 4226
rect 137006 4174 137058 4226
rect 139022 4174 139074 4226
rect 141262 4174 141314 4226
rect 141822 4174 141874 4226
rect 144958 4174 145010 4226
rect 146862 4174 146914 4226
rect 127598 4062 127650 4114
rect 19624 3894 19676 3946
rect 19728 3894 19780 3946
rect 19832 3894 19884 3946
rect 56444 3894 56496 3946
rect 56548 3894 56600 3946
rect 56652 3894 56704 3946
rect 93264 3894 93316 3946
rect 93368 3894 93420 3946
rect 93472 3894 93524 3946
rect 130084 3894 130136 3946
rect 130188 3894 130240 3946
rect 130292 3894 130344 3946
rect 8206 3614 8258 3666
rect 10222 3614 10274 3666
rect 11902 3614 11954 3666
rect 19966 3614 20018 3666
rect 21422 3614 21474 3666
rect 24558 3614 24610 3666
rect 28478 3614 28530 3666
rect 32398 3614 32450 3666
rect 36318 3614 36370 3666
rect 40238 3614 40290 3666
rect 43710 3614 43762 3666
rect 48078 3614 48130 3666
rect 51998 3614 52050 3666
rect 55470 3614 55522 3666
rect 59838 3614 59890 3666
rect 63758 3614 63810 3666
rect 67230 3614 67282 3666
rect 71374 3614 71426 3666
rect 72718 3614 72770 3666
rect 75518 3614 75570 3666
rect 76974 3614 77026 3666
rect 78766 3614 78818 3666
rect 80894 3614 80946 3666
rect 82686 3614 82738 3666
rect 86942 3614 86994 3666
rect 88734 3614 88786 3666
rect 90526 3614 90578 3666
rect 94110 3614 94162 3666
rect 97582 3614 97634 3666
rect 98590 3614 98642 3666
rect 99822 3614 99874 3666
rect 103742 3614 103794 3666
rect 105870 3614 105922 3666
rect 107662 3614 107714 3666
rect 109566 3614 109618 3666
rect 111806 3614 111858 3666
rect 116734 3614 116786 3666
rect 117630 3614 117682 3666
rect 119646 3614 119698 3666
rect 121550 3614 121602 3666
rect 123566 3614 123618 3666
rect 126478 3614 126530 3666
rect 128494 3614 128546 3666
rect 129278 3614 129330 3666
rect 129838 3614 129890 3666
rect 131182 3614 131234 3666
rect 133646 3614 133698 3666
rect 135102 3614 135154 3666
rect 139022 3614 139074 3666
rect 141486 3614 141538 3666
rect 143166 3614 143218 3666
rect 6974 3502 7026 3554
rect 8766 3502 8818 3554
rect 11006 3502 11058 3554
rect 12798 3502 12850 3554
rect 14926 3502 14978 3554
rect 16718 3502 16770 3554
rect 18734 3502 18786 3554
rect 20638 3502 20690 3554
rect 30270 3502 30322 3554
rect 73390 3502 73442 3554
rect 76302 3502 76354 3554
rect 78094 3502 78146 3554
rect 80222 3502 80274 3554
rect 82014 3502 82066 3554
rect 85374 3502 85426 3554
rect 86494 3502 86546 3554
rect 88174 3502 88226 3554
rect 89854 3502 89906 3554
rect 106318 3502 106370 3554
rect 106766 3502 106818 3554
rect 110350 3502 110402 3554
rect 113486 3502 113538 3554
rect 118078 3502 118130 3554
rect 133310 3502 133362 3554
rect 137006 3502 137058 3554
rect 137902 3502 137954 3554
rect 5854 3390 5906 3442
rect 13806 3390 13858 3442
rect 15598 3390 15650 3442
rect 17614 3390 17666 3442
rect 23438 3390 23490 3442
rect 25230 3390 25282 3442
rect 27134 3390 27186 3442
rect 29150 3390 29202 3442
rect 31390 3390 31442 3442
rect 33070 3390 33122 3442
rect 35198 3390 35250 3442
rect 36990 3390 37042 3442
rect 38894 3390 38946 3442
rect 40910 3390 40962 3442
rect 41918 3390 41970 3442
rect 42478 3390 42530 3442
rect 45390 3390 45442 3442
rect 46958 3390 47010 3442
rect 48750 3390 48802 3442
rect 50654 3390 50706 3442
rect 52670 3390 52722 3442
rect 53678 3390 53730 3442
rect 54238 3390 54290 3442
rect 57262 3390 57314 3442
rect 58718 3390 58770 3442
rect 60510 3390 60562 3442
rect 62414 3390 62466 3442
rect 64430 3390 64482 3442
rect 65438 3390 65490 3442
rect 65998 3390 66050 3442
rect 68910 3390 68962 3442
rect 70590 3390 70642 3442
rect 74510 3390 74562 3442
rect 84478 3390 84530 3442
rect 92318 3390 92370 3442
rect 92878 3390 92930 3442
rect 95230 3390 95282 3442
rect 96238 3390 96290 3442
rect 98030 3390 98082 3442
rect 99150 3390 99202 3442
rect 100830 3390 100882 3442
rect 103070 3390 103122 3442
rect 104750 3390 104802 3442
rect 108670 3390 108722 3442
rect 112590 3390 112642 3442
rect 113934 3390 113986 3442
rect 114830 3390 114882 3442
rect 115614 3390 115666 3442
rect 118526 3390 118578 3442
rect 120654 3390 120706 3442
rect 121998 3390 122050 3442
rect 122670 3390 122722 3442
rect 124350 3390 124402 3442
rect 126030 3390 126082 3442
rect 127374 3390 127426 3442
rect 130398 3390 130450 3442
rect 132190 3390 132242 3442
rect 134206 3390 134258 3442
rect 136110 3390 136162 3442
rect 140030 3390 140082 3442
rect 140926 3390 140978 3442
rect 141822 3390 141874 3442
rect 144174 3390 144226 3442
rect 145070 3390 145122 3442
rect 73166 3278 73218 3330
rect 86158 3278 86210 3330
rect 110686 3278 110738 3330
rect 138238 3278 138290 3330
rect 38034 3110 38086 3162
rect 38138 3110 38190 3162
rect 38242 3110 38294 3162
rect 74854 3110 74906 3162
rect 74958 3110 75010 3162
rect 75062 3110 75114 3162
rect 111674 3110 111726 3162
rect 111778 3110 111830 3162
rect 111882 3110 111934 3162
rect 148494 3110 148546 3162
rect 148598 3110 148650 3162
rect 148702 3110 148754 3162
<< metal2 >>
rect 147644 38836 147700 38846
rect 144508 37940 144564 37950
rect 19622 36876 19886 36886
rect 19678 36820 19726 36876
rect 19782 36820 19830 36876
rect 19622 36810 19886 36820
rect 56442 36876 56706 36886
rect 56498 36820 56546 36876
rect 56602 36820 56650 36876
rect 56442 36810 56706 36820
rect 93262 36876 93526 36886
rect 93318 36820 93366 36876
rect 93422 36820 93470 36876
rect 93262 36810 93526 36820
rect 130082 36876 130346 36886
rect 130138 36820 130186 36876
rect 130242 36820 130290 36876
rect 130082 36810 130346 36820
rect 144172 36596 144228 36606
rect 144508 36596 144564 37884
rect 144172 36594 144564 36596
rect 144172 36542 144174 36594
rect 144226 36542 144564 36594
rect 144172 36540 144564 36542
rect 144172 36530 144228 36540
rect 143052 36482 143108 36494
rect 143052 36430 143054 36482
rect 143106 36430 143108 36482
rect 139020 36260 139076 36270
rect 38032 36092 38296 36102
rect 38088 36036 38136 36092
rect 38192 36036 38240 36092
rect 38032 36026 38296 36036
rect 74852 36092 75116 36102
rect 74908 36036 74956 36092
rect 75012 36036 75060 36092
rect 74852 36026 75116 36036
rect 111672 36092 111936 36102
rect 111728 36036 111776 36092
rect 111832 36036 111880 36092
rect 111672 36026 111936 36036
rect 19622 35308 19886 35318
rect 19678 35252 19726 35308
rect 19782 35252 19830 35308
rect 19622 35242 19886 35252
rect 56442 35308 56706 35318
rect 56498 35252 56546 35308
rect 56602 35252 56650 35308
rect 56442 35242 56706 35252
rect 93262 35308 93526 35318
rect 93318 35252 93366 35308
rect 93422 35252 93470 35308
rect 93262 35242 93526 35252
rect 130082 35308 130346 35318
rect 130138 35252 130186 35308
rect 130242 35252 130290 35308
rect 130082 35242 130346 35252
rect 38032 34524 38296 34534
rect 38088 34468 38136 34524
rect 38192 34468 38240 34524
rect 38032 34458 38296 34468
rect 74852 34524 75116 34534
rect 74908 34468 74956 34524
rect 75012 34468 75060 34524
rect 74852 34458 75116 34468
rect 111672 34524 111936 34534
rect 111728 34468 111776 34524
rect 111832 34468 111880 34524
rect 111672 34458 111936 34468
rect 137340 34020 137396 34030
rect 19622 33740 19886 33750
rect 19678 33684 19726 33740
rect 19782 33684 19830 33740
rect 19622 33674 19886 33684
rect 56442 33740 56706 33750
rect 56498 33684 56546 33740
rect 56602 33684 56650 33740
rect 56442 33674 56706 33684
rect 93262 33740 93526 33750
rect 93318 33684 93366 33740
rect 93422 33684 93470 33740
rect 93262 33674 93526 33684
rect 130082 33740 130346 33750
rect 130138 33684 130186 33740
rect 130242 33684 130290 33740
rect 130082 33674 130346 33684
rect 134764 33124 134820 33134
rect 38032 32956 38296 32966
rect 38088 32900 38136 32956
rect 38192 32900 38240 32956
rect 38032 32890 38296 32900
rect 74852 32956 75116 32966
rect 74908 32900 74956 32956
rect 75012 32900 75060 32956
rect 74852 32890 75116 32900
rect 111672 32956 111936 32966
rect 111728 32900 111776 32956
rect 111832 32900 111880 32956
rect 111672 32890 111936 32900
rect 19622 32172 19886 32182
rect 19678 32116 19726 32172
rect 19782 32116 19830 32172
rect 19622 32106 19886 32116
rect 56442 32172 56706 32182
rect 56498 32116 56546 32172
rect 56602 32116 56650 32172
rect 56442 32106 56706 32116
rect 93262 32172 93526 32182
rect 93318 32116 93366 32172
rect 93422 32116 93470 32172
rect 93262 32106 93526 32116
rect 130082 32172 130346 32182
rect 130138 32116 130186 32172
rect 130242 32116 130290 32172
rect 130082 32106 130346 32116
rect 133308 31556 133364 31566
rect 38032 31388 38296 31398
rect 38088 31332 38136 31388
rect 38192 31332 38240 31388
rect 38032 31322 38296 31332
rect 74852 31388 75116 31398
rect 74908 31332 74956 31388
rect 75012 31332 75060 31388
rect 74852 31322 75116 31332
rect 111672 31388 111936 31398
rect 111728 31332 111776 31388
rect 111832 31332 111880 31388
rect 111672 31322 111936 31332
rect 131404 30884 131460 30894
rect 19622 30604 19886 30614
rect 19678 30548 19726 30604
rect 19782 30548 19830 30604
rect 19622 30538 19886 30548
rect 56442 30604 56706 30614
rect 56498 30548 56546 30604
rect 56602 30548 56650 30604
rect 56442 30538 56706 30548
rect 93262 30604 93526 30614
rect 93318 30548 93366 30604
rect 93422 30548 93470 30604
rect 93262 30538 93526 30548
rect 130082 30604 130346 30614
rect 130138 30548 130186 30604
rect 130242 30548 130290 30604
rect 130082 30538 130346 30548
rect 38032 29820 38296 29830
rect 38088 29764 38136 29820
rect 38192 29764 38240 29820
rect 38032 29754 38296 29764
rect 74852 29820 75116 29830
rect 74908 29764 74956 29820
rect 75012 29764 75060 29820
rect 74852 29754 75116 29764
rect 111672 29820 111936 29830
rect 111728 29764 111776 29820
rect 111832 29764 111880 29820
rect 111672 29754 111936 29764
rect 127932 29316 127988 29326
rect 19622 29036 19886 29046
rect 19678 28980 19726 29036
rect 19782 28980 19830 29036
rect 19622 28970 19886 28980
rect 56442 29036 56706 29046
rect 56498 28980 56546 29036
rect 56602 28980 56650 29036
rect 56442 28970 56706 28980
rect 93262 29036 93526 29046
rect 93318 28980 93366 29036
rect 93422 28980 93470 29036
rect 93262 28970 93526 28980
rect 38032 28252 38296 28262
rect 38088 28196 38136 28252
rect 38192 28196 38240 28252
rect 38032 28186 38296 28196
rect 74852 28252 75116 28262
rect 74908 28196 74956 28252
rect 75012 28196 75060 28252
rect 74852 28186 75116 28196
rect 111672 28252 111936 28262
rect 111728 28196 111776 28252
rect 111832 28196 111880 28252
rect 111672 28186 111936 28196
rect 124908 27748 124964 27758
rect 19622 27468 19886 27478
rect 19678 27412 19726 27468
rect 19782 27412 19830 27468
rect 19622 27402 19886 27412
rect 56442 27468 56706 27478
rect 56498 27412 56546 27468
rect 56602 27412 56650 27468
rect 56442 27402 56706 27412
rect 93262 27468 93526 27478
rect 93318 27412 93366 27468
rect 93422 27412 93470 27468
rect 93262 27402 93526 27412
rect 124124 26964 124180 26974
rect 38032 26684 38296 26694
rect 38088 26628 38136 26684
rect 38192 26628 38240 26684
rect 38032 26618 38296 26628
rect 74852 26684 75116 26694
rect 74908 26628 74956 26684
rect 75012 26628 75060 26684
rect 74852 26618 75116 26628
rect 111672 26684 111936 26694
rect 111728 26628 111776 26684
rect 111832 26628 111880 26684
rect 111672 26618 111936 26628
rect 19622 25900 19886 25910
rect 19678 25844 19726 25900
rect 19782 25844 19830 25900
rect 19622 25834 19886 25844
rect 56442 25900 56706 25910
rect 56498 25844 56546 25900
rect 56602 25844 56650 25900
rect 56442 25834 56706 25844
rect 93262 25900 93526 25910
rect 93318 25844 93366 25900
rect 93422 25844 93470 25900
rect 93262 25834 93526 25844
rect 120092 25172 120148 25182
rect 38032 25116 38296 25126
rect 38088 25060 38136 25116
rect 38192 25060 38240 25116
rect 38032 25050 38296 25060
rect 74852 25116 75116 25126
rect 74908 25060 74956 25116
rect 75012 25060 75060 25116
rect 74852 25050 75116 25060
rect 111672 25116 111936 25126
rect 111728 25060 111776 25116
rect 111832 25060 111880 25116
rect 111672 25050 111936 25060
rect 119196 24612 119252 24622
rect 19622 24332 19886 24342
rect 19678 24276 19726 24332
rect 19782 24276 19830 24332
rect 19622 24266 19886 24276
rect 56442 24332 56706 24342
rect 56498 24276 56546 24332
rect 56602 24276 56650 24332
rect 56442 24266 56706 24276
rect 93262 24332 93526 24342
rect 93318 24276 93366 24332
rect 93422 24276 93470 24332
rect 93262 24266 93526 24276
rect 38032 23548 38296 23558
rect 38088 23492 38136 23548
rect 38192 23492 38240 23548
rect 38032 23482 38296 23492
rect 74852 23548 75116 23558
rect 74908 23492 74956 23548
rect 75012 23492 75060 23548
rect 74852 23482 75116 23492
rect 111672 23548 111936 23558
rect 111728 23492 111776 23548
rect 111832 23492 111880 23548
rect 111672 23482 111936 23492
rect 19622 22764 19886 22774
rect 19678 22708 19726 22764
rect 19782 22708 19830 22764
rect 19622 22698 19886 22708
rect 56442 22764 56706 22774
rect 56498 22708 56546 22764
rect 56602 22708 56650 22764
rect 56442 22698 56706 22708
rect 93262 22764 93526 22774
rect 93318 22708 93366 22764
rect 93422 22708 93470 22764
rect 93262 22698 93526 22708
rect 113484 22148 113540 22158
rect 38032 21980 38296 21990
rect 38088 21924 38136 21980
rect 38192 21924 38240 21980
rect 38032 21914 38296 21924
rect 74852 21980 75116 21990
rect 74908 21924 74956 21980
rect 75012 21924 75060 21980
rect 74852 21914 75116 21924
rect 111672 21980 111936 21990
rect 111728 21924 111776 21980
rect 111832 21924 111880 21980
rect 111672 21914 111936 21924
rect 19622 21196 19886 21206
rect 19678 21140 19726 21196
rect 19782 21140 19830 21196
rect 19622 21130 19886 21140
rect 56442 21196 56706 21206
rect 56498 21140 56546 21196
rect 56602 21140 56650 21196
rect 56442 21130 56706 21140
rect 93262 21196 93526 21206
rect 93318 21140 93366 21196
rect 93422 21140 93470 21196
rect 93262 21130 93526 21140
rect 38032 20412 38296 20422
rect 38088 20356 38136 20412
rect 38192 20356 38240 20412
rect 38032 20346 38296 20356
rect 74852 20412 75116 20422
rect 74908 20356 74956 20412
rect 75012 20356 75060 20412
rect 74852 20346 75116 20356
rect 111672 20412 111936 20422
rect 111728 20356 111776 20412
rect 111832 20356 111880 20412
rect 111672 20346 111936 20356
rect 19622 19628 19886 19638
rect 19678 19572 19726 19628
rect 19782 19572 19830 19628
rect 19622 19562 19886 19572
rect 56442 19628 56706 19638
rect 56498 19572 56546 19628
rect 56602 19572 56650 19628
rect 56442 19562 56706 19572
rect 93262 19628 93526 19638
rect 93318 19572 93366 19628
rect 93422 19572 93470 19628
rect 93262 19562 93526 19572
rect 38032 18844 38296 18854
rect 38088 18788 38136 18844
rect 38192 18788 38240 18844
rect 38032 18778 38296 18788
rect 74852 18844 75116 18854
rect 74908 18788 74956 18844
rect 75012 18788 75060 18844
rect 74852 18778 75116 18788
rect 111672 18844 111936 18854
rect 111728 18788 111776 18844
rect 111832 18788 111880 18844
rect 111672 18778 111936 18788
rect 111580 18676 111636 18686
rect 111580 18582 111636 18620
rect 111244 18562 111300 18574
rect 111244 18510 111246 18562
rect 111298 18510 111300 18562
rect 110684 18338 110740 18350
rect 110684 18286 110686 18338
rect 110738 18286 110740 18338
rect 110684 18228 110740 18286
rect 111244 18228 111300 18510
rect 110684 18172 111300 18228
rect 19622 18060 19886 18070
rect 19678 18004 19726 18060
rect 19782 18004 19830 18060
rect 19622 17994 19886 18004
rect 56442 18060 56706 18070
rect 56498 18004 56546 18060
rect 56602 18004 56650 18060
rect 56442 17994 56706 18004
rect 93262 18060 93526 18070
rect 93318 18004 93366 18060
rect 93422 18004 93470 18060
rect 93262 17994 93526 18004
rect 106652 17444 106708 17454
rect 38032 17276 38296 17286
rect 38088 17220 38136 17276
rect 38192 17220 38240 17276
rect 38032 17210 38296 17220
rect 74852 17276 75116 17286
rect 74908 17220 74956 17276
rect 75012 17220 75060 17276
rect 74852 17210 75116 17220
rect 104524 16884 104580 16894
rect 19622 16492 19886 16502
rect 19678 16436 19726 16492
rect 19782 16436 19830 16492
rect 19622 16426 19886 16436
rect 56442 16492 56706 16502
rect 56498 16436 56546 16492
rect 56602 16436 56650 16492
rect 56442 16426 56706 16436
rect 93262 16492 93526 16502
rect 93318 16436 93366 16492
rect 93422 16436 93470 16492
rect 93262 16426 93526 16436
rect 103628 15876 103684 15886
rect 38032 15708 38296 15718
rect 38088 15652 38136 15708
rect 38192 15652 38240 15708
rect 38032 15642 38296 15652
rect 74852 15708 75116 15718
rect 74908 15652 74956 15708
rect 75012 15652 75060 15708
rect 74852 15642 75116 15652
rect 19622 14924 19886 14934
rect 19678 14868 19726 14924
rect 19782 14868 19830 14924
rect 19622 14858 19886 14868
rect 56442 14924 56706 14934
rect 56498 14868 56546 14924
rect 56602 14868 56650 14924
rect 56442 14858 56706 14868
rect 93262 14924 93526 14934
rect 93318 14868 93366 14924
rect 93422 14868 93470 14924
rect 93262 14858 93526 14868
rect 100492 14308 100548 14318
rect 38032 14140 38296 14150
rect 38088 14084 38136 14140
rect 38192 14084 38240 14140
rect 38032 14074 38296 14084
rect 74852 14140 75116 14150
rect 74908 14084 74956 14140
rect 75012 14084 75060 14140
rect 74852 14074 75116 14084
rect 19622 13356 19886 13366
rect 19678 13300 19726 13356
rect 19782 13300 19830 13356
rect 19622 13290 19886 13300
rect 56442 13356 56706 13366
rect 56498 13300 56546 13356
rect 56602 13300 56650 13356
rect 56442 13290 56706 13300
rect 93262 13356 93526 13366
rect 93318 13300 93366 13356
rect 93422 13300 93470 13356
rect 93262 13290 93526 13300
rect 100044 12852 100100 12862
rect 38032 12572 38296 12582
rect 38088 12516 38136 12572
rect 38192 12516 38240 12572
rect 38032 12506 38296 12516
rect 74852 12572 75116 12582
rect 74908 12516 74956 12572
rect 75012 12516 75060 12572
rect 74852 12506 75116 12516
rect 71372 12404 71428 12414
rect 63868 11956 63924 11966
rect 19622 11788 19886 11798
rect 19678 11732 19726 11788
rect 19782 11732 19830 11788
rect 19622 11722 19886 11732
rect 56442 11788 56706 11798
rect 56498 11732 56546 11788
rect 56602 11732 56650 11788
rect 56442 11722 56706 11732
rect 38032 11004 38296 11014
rect 38088 10948 38136 11004
rect 38192 10948 38240 11004
rect 38032 10938 38296 10948
rect 53900 10724 53956 10734
rect 32396 10612 32452 10622
rect 17052 10388 17108 10398
rect 12124 9044 12180 9054
rect 10780 7364 10836 7374
rect 9996 5124 10052 5134
rect 8764 4564 8820 4574
rect 8316 4340 8372 4350
rect 8316 4246 8372 4284
rect 6636 4228 6692 4238
rect 7196 4228 7252 4238
rect 6636 4226 7028 4228
rect 6636 4174 6638 4226
rect 6690 4174 7028 4226
rect 6636 4172 7028 4174
rect 6636 4162 6692 4172
rect 6972 3554 7028 4172
rect 6972 3502 6974 3554
rect 7026 3502 7028 3554
rect 5180 3444 5236 3454
rect 5180 800 5236 3388
rect 5852 3444 5908 3454
rect 5852 3350 5908 3388
rect 6972 3332 7028 3502
rect 6972 3266 7028 3276
rect 7084 4226 7252 4228
rect 7084 4174 7198 4226
rect 7250 4174 7252 4226
rect 7084 4172 7252 4174
rect 7084 980 7140 4172
rect 7196 4162 7252 4172
rect 8204 3668 8260 3678
rect 8204 3666 8596 3668
rect 8204 3614 8206 3666
rect 8258 3614 8596 3666
rect 8204 3612 8596 3614
rect 8204 3602 8260 3612
rect 6860 924 7140 980
rect 6860 800 6916 924
rect 8540 800 8596 3612
rect 8764 3554 8820 4508
rect 9772 4564 9828 4574
rect 9772 4470 9828 4508
rect 8876 4340 8932 4350
rect 8876 4246 8932 4284
rect 9996 4340 10052 5068
rect 10780 4564 10836 7308
rect 10780 4498 10836 4508
rect 11004 4564 11060 4574
rect 9996 4274 10052 4284
rect 8764 3502 8766 3554
rect 8818 3502 8820 3554
rect 8764 3490 8820 3502
rect 10220 3666 10276 3678
rect 10220 3614 10222 3666
rect 10274 3614 10276 3666
rect 10220 800 10276 3614
rect 11004 3554 11060 4508
rect 11340 4564 11396 4574
rect 11340 4470 11396 4508
rect 12124 4564 12180 8988
rect 15036 8932 15092 8942
rect 12124 4498 12180 4508
rect 13020 4564 13076 4574
rect 11004 3502 11006 3554
rect 11058 3502 11060 3554
rect 11004 3490 11060 3502
rect 11900 3666 11956 3678
rect 11900 3614 11902 3666
rect 11954 3614 11956 3666
rect 11900 800 11956 3614
rect 12796 3556 12852 3566
rect 13020 3556 13076 4508
rect 15036 4564 15092 8876
rect 15036 4498 15092 4508
rect 17052 4562 17108 10332
rect 19622 10220 19886 10230
rect 19678 10164 19726 10220
rect 19782 10164 19830 10220
rect 19622 10154 19886 10164
rect 19622 8652 19886 8662
rect 19678 8596 19726 8652
rect 19782 8596 19830 8652
rect 19622 8586 19886 8596
rect 19622 7084 19886 7094
rect 19678 7028 19726 7084
rect 19782 7028 19830 7084
rect 19622 7018 19886 7028
rect 30044 5908 30100 5918
rect 28588 5684 28644 5694
rect 19622 5516 19886 5526
rect 19678 5460 19726 5516
rect 19782 5460 19830 5516
rect 19622 5450 19886 5460
rect 17052 4510 17054 4562
rect 17106 4510 17108 4562
rect 15148 4226 15204 4238
rect 15148 4174 15150 4226
rect 15202 4174 15204 4226
rect 12796 3554 13076 3556
rect 12796 3502 12798 3554
rect 12850 3502 13076 3554
rect 12796 3500 13076 3502
rect 14924 3780 14980 3790
rect 14924 3554 14980 3724
rect 15148 3780 15204 4174
rect 15148 3714 15204 3724
rect 14924 3502 14926 3554
rect 14978 3502 14980 3554
rect 12796 3490 12852 3500
rect 14924 3490 14980 3502
rect 16716 3556 16772 3566
rect 17052 3556 17108 4510
rect 27132 5348 27188 5358
rect 22316 4452 22372 4462
rect 25788 4452 25844 4462
rect 21980 4450 22372 4452
rect 21980 4398 22318 4450
rect 22370 4398 22372 4450
rect 21980 4396 22372 4398
rect 20076 4338 20132 4350
rect 20076 4286 20078 4338
rect 20130 4286 20132 4338
rect 18284 4226 18340 4238
rect 18956 4228 19012 4238
rect 18284 4174 18286 4226
rect 18338 4174 18340 4226
rect 18284 3668 18340 4174
rect 18284 3602 18340 3612
rect 18620 4226 19012 4228
rect 18620 4174 18958 4226
rect 19010 4174 19012 4226
rect 18620 4172 19012 4174
rect 16716 3554 17108 3556
rect 16716 3502 16718 3554
rect 16770 3502 17108 3554
rect 16716 3500 17108 3502
rect 16716 3490 16772 3500
rect 13804 3444 13860 3454
rect 15596 3444 15652 3454
rect 13580 3442 13860 3444
rect 13580 3390 13806 3442
rect 13858 3390 13860 3442
rect 13580 3388 13860 3390
rect 13580 800 13636 3388
rect 13804 3378 13860 3388
rect 15260 3442 15652 3444
rect 15260 3390 15598 3442
rect 15650 3390 15652 3442
rect 15260 3388 15652 3390
rect 15260 800 15316 3388
rect 15596 3378 15652 3388
rect 17612 3442 17668 3454
rect 17612 3390 17614 3442
rect 17666 3390 17668 3442
rect 16940 924 17332 980
rect 16940 800 16996 924
rect 5152 0 5264 800
rect 6832 0 6944 800
rect 8512 0 8624 800
rect 10192 0 10304 800
rect 11872 0 11984 800
rect 13552 0 13664 800
rect 15232 0 15344 800
rect 16912 0 17024 800
rect 17276 756 17332 924
rect 17612 756 17668 3390
rect 18620 800 18676 4172
rect 18956 4162 19012 4172
rect 20076 4116 20132 4286
rect 20076 4050 20132 4060
rect 20524 4226 20580 4238
rect 20524 4174 20526 4226
rect 20578 4174 20580 4226
rect 20524 4116 20580 4174
rect 21756 4228 21812 4238
rect 21980 4228 22036 4396
rect 22316 4386 22372 4396
rect 25340 4450 25844 4452
rect 25340 4398 25790 4450
rect 25842 4398 25844 4450
rect 25340 4396 25844 4398
rect 21756 4226 22036 4228
rect 21756 4174 21758 4226
rect 21810 4174 22036 4226
rect 21756 4172 22036 4174
rect 21756 4162 21812 4172
rect 20524 4050 20580 4060
rect 19622 3948 19886 3958
rect 19678 3892 19726 3948
rect 19782 3892 19830 3948
rect 19622 3882 19886 3892
rect 20636 3892 20692 3902
rect 18732 3668 18788 3678
rect 18732 3554 18788 3612
rect 19964 3668 20020 3678
rect 19964 3666 20356 3668
rect 19964 3614 19966 3666
rect 20018 3614 20356 3666
rect 19964 3612 20356 3614
rect 19964 3602 20020 3612
rect 18732 3502 18734 3554
rect 18786 3502 18788 3554
rect 18732 3490 18788 3502
rect 20300 800 20356 3612
rect 20636 3554 20692 3836
rect 21420 3892 21476 3902
rect 21420 3666 21476 3836
rect 21420 3614 21422 3666
rect 21474 3614 21476 3666
rect 21420 3602 21476 3614
rect 20636 3502 20638 3554
rect 20690 3502 20692 3554
rect 20636 3490 20692 3502
rect 21980 800 22036 4172
rect 23660 4228 23716 4238
rect 25004 4228 25060 4238
rect 25340 4228 25396 4396
rect 25788 4386 25844 4396
rect 23660 4226 23828 4228
rect 23660 4174 23662 4226
rect 23714 4174 23828 4226
rect 23660 4172 23828 4174
rect 23660 4162 23716 4172
rect 23436 3444 23492 3454
rect 23660 3444 23716 3454
rect 23436 3442 23660 3444
rect 23436 3390 23438 3442
rect 23490 3390 23660 3442
rect 23436 3388 23660 3390
rect 23436 3378 23492 3388
rect 23660 800 23716 3388
rect 23772 2436 23828 4172
rect 25004 4226 25396 4228
rect 25004 4174 25006 4226
rect 25058 4174 25396 4226
rect 25004 4172 25396 4174
rect 25004 4162 25060 4172
rect 23772 2370 23828 2380
rect 24556 3666 24612 3678
rect 24556 3614 24558 3666
rect 24610 3614 24612 3666
rect 24556 1652 24612 3614
rect 25228 3444 25284 3454
rect 25228 3350 25284 3388
rect 24556 1586 24612 1596
rect 25340 800 25396 4172
rect 27132 4226 27188 5292
rect 27132 4174 27134 4226
rect 27186 4174 27188 4226
rect 27132 4162 27188 4174
rect 28476 3668 28532 3678
rect 28588 3668 28644 5628
rect 28476 3666 28644 3668
rect 28476 3614 28478 3666
rect 28530 3614 28644 3666
rect 28476 3612 28644 3614
rect 28700 4450 28756 4462
rect 28700 4398 28702 4450
rect 28754 4398 28756 4450
rect 28476 3602 28532 3612
rect 28700 3556 28756 4398
rect 30044 4226 30100 5852
rect 30044 4174 30046 4226
rect 30098 4174 30100 4226
rect 30044 4162 30100 4174
rect 30380 4898 30436 4910
rect 30380 4846 30382 4898
rect 30434 4846 30436 4898
rect 30380 4452 30436 4846
rect 30716 4452 30772 4462
rect 30380 4450 30772 4452
rect 30380 4398 30718 4450
rect 30770 4398 30772 4450
rect 30380 4396 30772 4398
rect 27132 3444 27188 3454
rect 27020 3388 27132 3444
rect 27020 800 27076 3388
rect 27132 3312 27188 3388
rect 28700 800 28756 3500
rect 30268 3556 30324 3566
rect 30268 3462 30324 3500
rect 29148 3444 29204 3454
rect 29148 3350 29204 3388
rect 30380 800 30436 4396
rect 30716 4386 30772 4396
rect 31948 4226 32004 4238
rect 31948 4174 31950 4226
rect 32002 4174 32004 4226
rect 31388 3444 31444 3454
rect 31388 3350 31444 3388
rect 31948 2324 32004 4174
rect 32396 3666 32452 10556
rect 38032 9436 38296 9446
rect 38088 9380 38136 9436
rect 38192 9380 38240 9436
rect 38032 9370 38296 9380
rect 47180 9156 47236 9166
rect 38032 7868 38296 7878
rect 38088 7812 38136 7868
rect 38192 7812 38240 7868
rect 38032 7802 38296 7812
rect 36316 7252 36372 7262
rect 34076 4452 34132 4462
rect 33740 4450 34132 4452
rect 33740 4398 34078 4450
rect 34130 4398 34132 4450
rect 33740 4396 34132 4398
rect 32956 4228 33012 4238
rect 32956 4134 33012 4172
rect 33740 4228 33796 4396
rect 34076 4386 34132 4396
rect 32396 3614 32398 3666
rect 32450 3614 32452 3666
rect 32396 3602 32452 3614
rect 31948 2258 32004 2268
rect 32060 3444 32116 3454
rect 32060 800 32116 3388
rect 33068 3444 33124 3454
rect 33068 3350 33124 3388
rect 33740 800 33796 4172
rect 35420 4228 35476 4238
rect 35420 4226 35700 4228
rect 35420 4174 35422 4226
rect 35474 4174 35700 4226
rect 35420 4172 35700 4174
rect 35420 4162 35476 4172
rect 35196 3444 35252 3454
rect 35420 3444 35476 3454
rect 35196 3442 35420 3444
rect 35196 3390 35198 3442
rect 35250 3390 35420 3442
rect 35196 3388 35420 3390
rect 35196 3378 35252 3388
rect 35420 800 35476 3388
rect 35644 868 35700 4172
rect 36316 3666 36372 7196
rect 40348 6804 40404 6814
rect 38032 6300 38296 6310
rect 38088 6244 38136 6300
rect 38192 6244 38240 6300
rect 38032 6234 38296 6244
rect 38032 4732 38296 4742
rect 38088 4676 38136 4732
rect 38192 4676 38240 4732
rect 38032 4666 38296 4676
rect 37436 4452 37492 4462
rect 37100 4450 37492 4452
rect 37100 4398 37438 4450
rect 37490 4398 37492 4450
rect 37100 4396 37492 4398
rect 36876 4228 36932 4238
rect 37100 4228 37156 4396
rect 37436 4386 37492 4396
rect 36876 4226 37156 4228
rect 36876 4174 36878 4226
rect 36930 4174 37156 4226
rect 36876 4172 37156 4174
rect 36876 4162 36932 4172
rect 36316 3614 36318 3666
rect 36370 3614 36372 3666
rect 36316 3602 36372 3614
rect 36988 3444 37044 3454
rect 36988 3350 37044 3388
rect 35644 802 35700 812
rect 37100 800 37156 4172
rect 38668 4226 38724 4238
rect 38668 4174 38670 4226
rect 38722 4174 38724 4226
rect 38032 3164 38296 3174
rect 38088 3108 38136 3164
rect 38192 3108 38240 3164
rect 38032 3098 38296 3108
rect 38668 2660 38724 4174
rect 40236 3668 40292 3678
rect 40348 3668 40404 6748
rect 45500 4898 45556 4910
rect 45500 4846 45502 4898
rect 45554 4846 45556 4898
rect 40796 4452 40852 4462
rect 40796 4228 40852 4396
rect 41692 4452 41748 4462
rect 41692 4358 41748 4396
rect 43820 4450 43876 4462
rect 43820 4398 43822 4450
rect 43874 4398 43876 4450
rect 40236 3666 40404 3668
rect 40236 3614 40238 3666
rect 40290 3614 40404 3666
rect 40236 3612 40404 3614
rect 40460 4226 40852 4228
rect 40460 4174 40798 4226
rect 40850 4174 40852 4226
rect 40460 4172 40852 4174
rect 40236 3602 40292 3612
rect 38892 3444 38948 3454
rect 38668 2594 38724 2604
rect 38780 3388 38892 3444
rect 38780 800 38836 3388
rect 38892 3312 38948 3388
rect 40460 800 40516 4172
rect 40796 4162 40852 4172
rect 43036 4226 43092 4238
rect 43036 4174 43038 4226
rect 43090 4174 43092 4226
rect 40908 3444 40964 3454
rect 40908 3350 40964 3388
rect 41916 3444 41972 3454
rect 42476 3444 42532 3454
rect 41916 3442 42532 3444
rect 41916 3390 41918 3442
rect 41970 3390 42478 3442
rect 42530 3390 42532 3442
rect 41916 3388 42532 3390
rect 41916 3378 41972 3388
rect 42140 800 42196 3388
rect 42476 3378 42532 3388
rect 43036 2884 43092 4174
rect 43036 2818 43092 2828
rect 43708 3666 43764 3678
rect 43708 3614 43710 3666
rect 43762 3614 43764 3666
rect 43708 1092 43764 3614
rect 43708 1026 43764 1036
rect 43820 3444 43876 4398
rect 45500 4452 45556 4846
rect 45836 4452 45892 4462
rect 45500 4450 45892 4452
rect 45500 4398 45838 4450
rect 45890 4398 45892 4450
rect 45500 4396 45892 4398
rect 43820 800 43876 3388
rect 45164 4226 45220 4238
rect 45164 4174 45166 4226
rect 45218 4174 45220 4226
rect 45164 1540 45220 4174
rect 45388 3444 45444 3454
rect 45388 3350 45444 3388
rect 45164 1474 45220 1484
rect 45500 800 45556 4396
rect 45836 4386 45892 4396
rect 47180 4226 47236 9100
rect 50988 7588 51044 7598
rect 47180 4174 47182 4226
rect 47234 4174 47236 4226
rect 47180 4162 47236 4174
rect 48860 4452 48916 4462
rect 48860 4226 48916 4396
rect 49644 4452 49700 4462
rect 49644 4358 49700 4396
rect 48860 4174 48862 4226
rect 48914 4174 48916 4226
rect 48076 3666 48132 3678
rect 48076 3614 48078 3666
rect 48130 3614 48132 3666
rect 46956 3444 47012 3454
rect 47180 3444 47236 3454
rect 46956 3442 47180 3444
rect 46956 3390 46958 3442
rect 47010 3390 47180 3442
rect 46956 3388 47180 3390
rect 46956 3378 47012 3388
rect 47180 800 47236 3388
rect 48076 2772 48132 3614
rect 48748 3444 48804 3454
rect 48748 3350 48804 3388
rect 48076 2706 48132 2716
rect 48860 800 48916 4174
rect 50988 4226 51044 7532
rect 52556 4452 52612 4462
rect 52220 4450 52612 4452
rect 52220 4398 52558 4450
rect 52610 4398 52612 4450
rect 52220 4396 52612 4398
rect 50988 4174 50990 4226
rect 51042 4174 51044 4226
rect 50988 4162 51044 4174
rect 51996 4228 52052 4238
rect 52220 4228 52276 4396
rect 52556 4386 52612 4396
rect 51996 4226 52276 4228
rect 51996 4174 51998 4226
rect 52050 4174 52276 4226
rect 51996 4172 52276 4174
rect 51996 4162 52052 4172
rect 51996 3668 52052 3678
rect 51996 3666 52164 3668
rect 51996 3614 51998 3666
rect 52050 3614 52164 3666
rect 51996 3612 52164 3614
rect 51996 3602 52052 3612
rect 50652 3444 50708 3454
rect 50540 3388 50652 3444
rect 50540 800 50596 3388
rect 50652 3312 50708 3388
rect 52108 1316 52164 3612
rect 52108 1250 52164 1260
rect 52220 800 52276 4172
rect 53900 4226 53956 10668
rect 56442 10220 56706 10230
rect 56498 10164 56546 10220
rect 56602 10164 56650 10220
rect 56442 10154 56706 10164
rect 56442 8652 56706 8662
rect 56498 8596 56546 8652
rect 56602 8596 56650 8652
rect 56442 8586 56706 8596
rect 57036 8484 57092 8494
rect 56442 7084 56706 7094
rect 56498 7028 56546 7084
rect 56602 7028 56650 7084
rect 56442 7018 56706 7028
rect 56442 5516 56706 5526
rect 56498 5460 56546 5516
rect 56602 5460 56650 5516
rect 56442 5450 56706 5460
rect 56924 4898 56980 4910
rect 56924 4846 56926 4898
rect 56978 4846 56980 4898
rect 53900 4174 53902 4226
rect 53954 4174 53956 4226
rect 53900 4162 53956 4174
rect 55580 4452 55636 4462
rect 56924 4452 56980 4846
rect 55580 4450 56980 4452
rect 55580 4398 55582 4450
rect 55634 4398 56980 4450
rect 55580 4396 56980 4398
rect 55468 3666 55524 3678
rect 55468 3614 55470 3666
rect 55522 3614 55524 3666
rect 52668 3444 52724 3454
rect 52668 3350 52724 3388
rect 53676 3444 53732 3454
rect 54236 3444 54292 3454
rect 53676 3442 54292 3444
rect 53676 3390 53678 3442
rect 53730 3390 54238 3442
rect 54290 3390 54292 3442
rect 53676 3388 54292 3390
rect 53676 3378 53732 3388
rect 53900 800 53956 3388
rect 54236 3378 54292 3388
rect 55468 2996 55524 3614
rect 55468 2930 55524 2940
rect 55580 800 55636 4396
rect 56700 4228 56756 4238
rect 57036 4228 57092 8428
rect 59836 6916 59892 6926
rect 57596 4452 57652 4462
rect 56700 4226 57092 4228
rect 56700 4174 56702 4226
rect 56754 4174 57092 4226
rect 56700 4172 57092 4174
rect 57260 4450 57652 4452
rect 57260 4398 57598 4450
rect 57650 4398 57652 4450
rect 57260 4396 57652 4398
rect 56700 4162 56756 4172
rect 56442 3948 56706 3958
rect 56498 3892 56546 3948
rect 56602 3892 56650 3948
rect 56442 3882 56706 3892
rect 57260 3442 57316 4396
rect 57596 4386 57652 4396
rect 58940 4228 58996 4238
rect 58940 4226 59108 4228
rect 58940 4174 58942 4226
rect 58994 4174 59108 4226
rect 58940 4172 59108 4174
rect 58940 4162 58996 4172
rect 57260 3390 57262 3442
rect 57314 3390 57316 3442
rect 57260 800 57316 3390
rect 58716 3444 58772 3454
rect 58940 3444 58996 3454
rect 58716 3442 58940 3444
rect 58716 3390 58718 3442
rect 58770 3390 58940 3442
rect 58716 3388 58940 3390
rect 58716 3378 58772 3388
rect 58940 800 58996 3388
rect 59052 1204 59108 4172
rect 59836 3666 59892 6860
rect 63756 5122 63812 5134
rect 63756 5070 63758 5122
rect 63810 5070 63812 5122
rect 63756 4900 63812 5070
rect 63756 4834 63812 4844
rect 60956 4452 61012 4462
rect 60620 4450 61012 4452
rect 60620 4398 60958 4450
rect 61010 4398 61012 4450
rect 60620 4396 61012 4398
rect 60396 4228 60452 4238
rect 60620 4228 60676 4396
rect 60956 4386 61012 4396
rect 60396 4226 60676 4228
rect 60396 4174 60398 4226
rect 60450 4174 60676 4226
rect 60396 4172 60676 4174
rect 60396 4162 60452 4172
rect 59836 3614 59838 3666
rect 59890 3614 59892 3666
rect 59836 3602 59892 3614
rect 60508 3444 60564 3454
rect 60508 3350 60564 3388
rect 59052 1138 59108 1148
rect 60620 800 60676 4172
rect 62188 4226 62244 4238
rect 62188 4174 62190 4226
rect 62242 4174 62244 4226
rect 62188 2548 62244 4174
rect 63756 3668 63812 3678
rect 63868 3668 63924 11900
rect 70588 6020 70644 6030
rect 65660 5236 65716 5246
rect 65660 5142 65716 5180
rect 64316 5010 64372 5022
rect 64316 4958 64318 5010
rect 64370 4958 64372 5010
rect 63756 3666 63924 3668
rect 63756 3614 63758 3666
rect 63810 3614 63924 3666
rect 63756 3612 63924 3614
rect 63980 4900 64036 4910
rect 63756 3602 63812 3612
rect 62412 3444 62468 3454
rect 62188 2482 62244 2492
rect 62300 3388 62412 3444
rect 62300 800 62356 3388
rect 62412 3312 62468 3388
rect 63980 800 64036 4844
rect 64316 4900 64372 4958
rect 64316 4834 64372 4844
rect 69356 4898 69412 4910
rect 69356 4846 69358 4898
rect 69410 4846 69412 4898
rect 64092 4564 64148 4574
rect 64092 2660 64148 4508
rect 67340 4450 67396 4462
rect 69356 4452 69412 4846
rect 67340 4398 67342 4450
rect 67394 4398 67396 4450
rect 67228 3666 67284 3678
rect 67228 3614 67230 3666
rect 67282 3614 67284 3666
rect 64428 3444 64484 3454
rect 64428 3350 64484 3388
rect 65436 3444 65492 3454
rect 65996 3444 66052 3454
rect 65436 3442 66052 3444
rect 65436 3390 65438 3442
rect 65490 3390 65998 3442
rect 66050 3390 66052 3442
rect 65436 3388 66052 3390
rect 65436 3378 65492 3388
rect 64092 2594 64148 2604
rect 65660 800 65716 3388
rect 65996 3378 66052 3388
rect 67228 980 67284 3614
rect 67228 914 67284 924
rect 67340 3444 67396 4398
rect 69020 4450 69412 4452
rect 69020 4398 69358 4450
rect 69410 4398 69412 4450
rect 69020 4396 69412 4398
rect 67340 800 67396 3388
rect 68684 4226 68740 4238
rect 68684 4174 68686 4226
rect 68738 4174 68740 4226
rect 68684 1428 68740 4174
rect 68908 3444 68964 3454
rect 68908 3350 68964 3388
rect 68684 1362 68740 1372
rect 69020 800 69076 4396
rect 69356 4386 69412 4396
rect 70588 4226 70644 5964
rect 70588 4174 70590 4226
rect 70642 4174 70644 4226
rect 70588 4162 70644 4174
rect 70700 4228 70756 4238
rect 70588 3444 70644 3454
rect 70700 3444 70756 4172
rect 71372 3666 71428 12348
rect 82796 12292 82852 12302
rect 74852 11004 75116 11014
rect 74908 10948 74956 11004
rect 75012 10948 75060 11004
rect 74852 10938 75116 10948
rect 74732 10500 74788 10510
rect 74508 5796 74564 5806
rect 73836 5124 73892 5134
rect 73388 5012 73444 5022
rect 72604 4452 72660 4462
rect 71820 4228 71876 4238
rect 72604 4228 72660 4396
rect 71820 4134 71876 4172
rect 72380 4226 72660 4228
rect 72380 4174 72606 4226
rect 72658 4174 72660 4226
rect 72380 4172 72660 4174
rect 71372 3614 71374 3666
rect 71426 3614 71428 3666
rect 71372 3602 71428 3614
rect 70588 3442 70756 3444
rect 70588 3390 70590 3442
rect 70642 3390 70756 3442
rect 70588 3388 70756 3390
rect 70588 3378 70644 3388
rect 70700 800 70756 3388
rect 72380 800 72436 4172
rect 72604 4162 72660 4172
rect 72716 3892 72772 3902
rect 72716 3666 72772 3836
rect 72716 3614 72718 3666
rect 72770 3614 72772 3666
rect 72716 3602 72772 3614
rect 73388 3892 73444 4956
rect 73500 4452 73556 4462
rect 73500 4358 73556 4396
rect 73836 4452 73892 5068
rect 73836 4386 73892 4396
rect 73388 3554 73444 3836
rect 73388 3502 73390 3554
rect 73442 3502 73444 3554
rect 73388 3490 73444 3502
rect 74508 3444 74564 5740
rect 74732 4226 74788 10444
rect 79436 9604 79492 9614
rect 74852 9436 75116 9446
rect 74908 9380 74956 9436
rect 75012 9380 75060 9436
rect 74852 9370 75116 9380
rect 75628 8820 75684 8830
rect 74852 7868 75116 7878
rect 74908 7812 74956 7868
rect 75012 7812 75060 7868
rect 74852 7802 75116 7812
rect 74852 6300 75116 6310
rect 74908 6244 74956 6300
rect 75012 6244 75060 6300
rect 74852 6234 75116 6244
rect 75404 5012 75460 5022
rect 75404 4918 75460 4956
rect 74852 4732 75116 4742
rect 74908 4676 74956 4732
rect 75012 4676 75060 4732
rect 74852 4666 75116 4676
rect 75628 4676 75684 8764
rect 76188 8036 76244 8046
rect 75740 5796 75796 5806
rect 75740 5702 75796 5740
rect 76188 5234 76244 7980
rect 77980 7364 78036 7374
rect 76188 5182 76190 5234
rect 76242 5182 76244 5234
rect 76188 5012 76244 5182
rect 76188 4946 76244 4956
rect 77196 5460 77252 5470
rect 75740 4900 75796 4910
rect 75740 4898 75908 4900
rect 75740 4846 75742 4898
rect 75794 4846 75908 4898
rect 75740 4844 75908 4846
rect 75740 4834 75796 4844
rect 75628 4620 75796 4676
rect 75628 4452 75684 4462
rect 75628 4358 75684 4396
rect 74732 4174 74734 4226
rect 74786 4174 74788 4226
rect 74732 4162 74788 4174
rect 75740 3892 75796 4620
rect 75628 3836 75796 3892
rect 75516 3668 75572 3678
rect 75628 3668 75684 3836
rect 75516 3666 75684 3668
rect 75516 3614 75518 3666
rect 75570 3614 75684 3666
rect 75516 3612 75684 3614
rect 75740 3668 75796 3678
rect 75516 3602 75572 3612
rect 74060 3442 74564 3444
rect 74060 3390 74510 3442
rect 74562 3390 74564 3442
rect 74060 3388 74564 3390
rect 73164 3332 73220 3342
rect 73164 3238 73220 3276
rect 74060 800 74116 3388
rect 74508 3378 74564 3388
rect 74852 3164 75116 3174
rect 74908 3108 74956 3164
rect 75012 3108 75060 3164
rect 74852 3098 75116 3108
rect 75740 800 75796 3612
rect 75852 3556 75908 4844
rect 76524 4564 76580 4574
rect 77196 4564 77252 5404
rect 77644 5460 77700 5470
rect 77644 5234 77700 5404
rect 77644 5182 77646 5234
rect 77698 5182 77700 5234
rect 77644 5170 77700 5182
rect 75964 4562 77252 4564
rect 75964 4510 76526 4562
rect 76578 4510 77252 4562
rect 75964 4508 77252 4510
rect 75964 4450 76020 4508
rect 76524 4498 76580 4508
rect 75964 4398 75966 4450
rect 76018 4398 76020 4450
rect 75964 4386 76020 4398
rect 77196 4338 77252 4508
rect 77980 4562 78036 7308
rect 79436 5234 79492 9548
rect 79436 5182 79438 5234
rect 79490 5182 79492 5234
rect 78540 5124 78596 5134
rect 77980 4510 77982 4562
rect 78034 4510 78036 4562
rect 77980 4498 78036 4510
rect 78316 5068 78540 5124
rect 77420 4452 77476 4462
rect 77420 4450 77588 4452
rect 77420 4398 77422 4450
rect 77474 4398 77588 4450
rect 77420 4396 77588 4398
rect 77420 4386 77476 4396
rect 77196 4286 77198 4338
rect 77250 4286 77252 4338
rect 77196 4274 77252 4286
rect 76972 3668 77028 3678
rect 76972 3574 77028 3612
rect 77420 3668 77476 3678
rect 76300 3556 76356 3566
rect 75852 3554 76356 3556
rect 75852 3502 76302 3554
rect 76354 3502 76356 3554
rect 75852 3500 76356 3502
rect 76300 3490 76356 3500
rect 77420 800 77476 3612
rect 77532 3556 77588 4396
rect 78316 4450 78372 5068
rect 78540 5030 78596 5068
rect 78876 5124 78932 5134
rect 78316 4398 78318 4450
rect 78370 4398 78372 4450
rect 78316 4386 78372 4398
rect 78876 4450 78932 5068
rect 79436 5124 79492 5182
rect 79436 5058 79492 5068
rect 79772 9044 79828 9054
rect 79772 4562 79828 8988
rect 80668 8932 80724 8942
rect 80556 7476 80612 7486
rect 80556 5460 80612 7420
rect 80556 5394 80612 5404
rect 80668 5010 80724 8876
rect 82796 6130 82852 12236
rect 98476 12180 98532 12190
rect 93262 11788 93526 11798
rect 93318 11732 93366 11788
rect 93422 11732 93470 11788
rect 93262 11722 93526 11732
rect 98028 11172 98084 11182
rect 85596 10388 85652 10398
rect 82796 6078 82798 6130
rect 82850 6078 82852 6130
rect 81004 5124 81060 5134
rect 81004 5030 81060 5068
rect 81452 5124 81508 5134
rect 81452 5030 81508 5068
rect 82236 5124 82292 5134
rect 82236 5030 82292 5068
rect 82796 5124 82852 6078
rect 85372 6244 85428 6254
rect 82796 5058 82852 5068
rect 83356 5124 83412 5134
rect 83356 5030 83412 5068
rect 83804 5124 83860 5134
rect 83804 5030 83860 5068
rect 84588 5124 84644 5134
rect 80668 4958 80670 5010
rect 80722 4958 80724 5010
rect 80668 4946 80724 4958
rect 79772 4510 79774 4562
rect 79826 4510 79828 4562
rect 79772 4498 79828 4510
rect 82460 4898 82516 4910
rect 82460 4846 82462 4898
rect 82514 4846 82516 4898
rect 78876 4398 78878 4450
rect 78930 4398 78932 4450
rect 78876 4386 78932 4398
rect 79212 4450 79268 4462
rect 79212 4398 79214 4450
rect 79266 4398 79268 4450
rect 78988 4228 79044 4238
rect 78988 3780 79044 4172
rect 78988 3714 79044 3724
rect 78764 3668 78820 3678
rect 78764 3574 78820 3612
rect 79100 3668 79156 3678
rect 78092 3556 78148 3566
rect 77532 3554 78148 3556
rect 77532 3502 78094 3554
rect 78146 3502 78148 3554
rect 77532 3500 78148 3502
rect 78092 3490 78148 3500
rect 79100 800 79156 3612
rect 79212 3556 79268 4398
rect 81676 4450 81732 4462
rect 81676 4398 81678 4450
rect 81730 4398 81732 4450
rect 80108 4340 80164 4350
rect 80108 4246 80164 4284
rect 80556 4340 80612 4350
rect 80556 4246 80612 4284
rect 81452 4340 81508 4350
rect 81452 4246 81508 4284
rect 80780 4004 80836 4014
rect 80220 3556 80276 3566
rect 79212 3554 80276 3556
rect 79212 3502 80222 3554
rect 80274 3502 80276 3554
rect 79212 3500 80276 3502
rect 80220 3490 80276 3500
rect 80780 800 80836 3948
rect 80892 3668 80948 3678
rect 80892 3574 80948 3612
rect 81676 3556 81732 4398
rect 82124 4340 82180 4350
rect 82460 4340 82516 4846
rect 83020 4898 83076 4910
rect 83020 4846 83022 4898
rect 83074 4846 83076 4898
rect 82684 4340 82740 4350
rect 82460 4338 82740 4340
rect 82460 4286 82686 4338
rect 82738 4286 82740 4338
rect 82460 4284 82740 4286
rect 82124 4226 82180 4284
rect 82684 4274 82740 4284
rect 82124 4174 82126 4226
rect 82178 4174 82180 4226
rect 82012 3556 82068 3566
rect 81676 3554 82068 3556
rect 81676 3502 82014 3554
rect 82066 3502 82068 3554
rect 81676 3500 82068 3502
rect 82012 3490 82068 3500
rect 82124 2660 82180 4174
rect 83020 4228 83076 4846
rect 83916 4900 83972 4910
rect 83020 4162 83076 4172
rect 83356 4226 83412 4238
rect 83356 4174 83358 4226
rect 83410 4174 83412 4226
rect 82684 4004 82740 4014
rect 82684 3666 82740 3948
rect 82684 3614 82686 3666
rect 82738 3614 82740 3666
rect 82684 3602 82740 3614
rect 82124 2594 82180 2604
rect 82460 3444 82516 3454
rect 82460 800 82516 3388
rect 83356 3444 83412 4174
rect 83356 3378 83412 3388
rect 83916 868 83972 4844
rect 84588 4338 84644 5068
rect 85372 5124 85428 6188
rect 85372 4562 85428 5068
rect 85484 5012 85540 5022
rect 85484 4918 85540 4956
rect 85372 4510 85374 4562
rect 85426 4510 85428 4562
rect 85372 4498 85428 4510
rect 84588 4286 84590 4338
rect 84642 4286 84644 4338
rect 84588 4274 84644 4286
rect 84812 4450 84868 4462
rect 84812 4398 84814 4450
rect 84866 4398 84868 4450
rect 84812 3556 84868 4398
rect 85372 3556 85428 3566
rect 84812 3554 85428 3556
rect 84812 3502 85374 3554
rect 85426 3502 85428 3554
rect 84812 3500 85428 3502
rect 85372 3490 85428 3500
rect 84476 3444 84532 3454
rect 83916 802 83972 812
rect 84140 3442 84532 3444
rect 84140 3390 84478 3442
rect 84530 3390 84532 3442
rect 84140 3388 84532 3390
rect 84140 800 84196 3388
rect 84476 3378 84532 3388
rect 85596 3332 85652 10332
rect 87164 10388 87220 10398
rect 86940 6132 86996 6142
rect 86716 6076 86940 6132
rect 86044 5796 86100 5806
rect 86044 5012 86100 5740
rect 86716 5122 86772 6076
rect 86940 6038 86996 6076
rect 86716 5070 86718 5122
rect 86770 5070 86772 5122
rect 86716 5058 86772 5070
rect 86940 5796 86996 5806
rect 86044 4946 86100 4956
rect 85820 4898 85876 4910
rect 85820 4846 85822 4898
rect 85874 4846 85876 4898
rect 85820 4340 85876 4846
rect 86380 4898 86436 4910
rect 86380 4846 86382 4898
rect 86434 4846 86436 4898
rect 86044 4340 86100 4350
rect 85820 4338 86100 4340
rect 85820 4286 86046 4338
rect 86098 4286 86100 4338
rect 85820 4284 86100 4286
rect 86044 4274 86100 4284
rect 86380 4004 86436 4846
rect 86380 3938 86436 3948
rect 86716 4226 86772 4238
rect 86716 4174 86718 4226
rect 86770 4174 86772 4226
rect 85596 3266 85652 3276
rect 85820 3892 85876 3902
rect 85820 800 85876 3836
rect 86716 3892 86772 4174
rect 86716 3826 86772 3836
rect 86940 3668 86996 5740
rect 87164 5236 87220 10332
rect 93262 10220 93526 10230
rect 93318 10164 93366 10220
rect 93422 10164 93470 10220
rect 93262 10154 93526 10164
rect 90748 9940 90804 9950
rect 90300 8932 90356 8942
rect 88396 6692 88452 6702
rect 87164 5170 87220 5180
rect 87836 6132 87892 6142
rect 87724 5012 87780 5022
rect 87724 4918 87780 4956
rect 87388 4898 87444 4910
rect 87388 4846 87390 4898
rect 87442 4846 87444 4898
rect 87388 4116 87444 4846
rect 87836 4450 87892 6076
rect 88396 6132 88452 6636
rect 88396 6000 88452 6076
rect 88956 5908 89012 5918
rect 88172 5012 88228 5022
rect 88172 4900 88228 4956
rect 88956 5012 89012 5852
rect 89404 5236 89460 5246
rect 89404 5122 89460 5180
rect 89852 5236 89908 5246
rect 89852 5142 89908 5180
rect 90188 5236 90244 5246
rect 89404 5070 89406 5122
rect 89458 5070 89460 5122
rect 89404 5058 89460 5070
rect 88956 4946 89012 4956
rect 88172 4898 88340 4900
rect 88172 4846 88174 4898
rect 88226 4846 88340 4898
rect 88172 4844 88340 4846
rect 88172 4834 88228 4844
rect 87836 4398 87838 4450
rect 87890 4398 87892 4450
rect 87836 4386 87892 4398
rect 88172 4450 88228 4462
rect 88172 4398 88174 4450
rect 88226 4398 88228 4450
rect 87388 4050 87444 4060
rect 86492 3666 86996 3668
rect 86492 3614 86942 3666
rect 86994 3614 86996 3666
rect 86492 3612 86996 3614
rect 86492 3554 86548 3612
rect 86940 3602 86996 3612
rect 87500 3668 87556 3678
rect 86492 3502 86494 3554
rect 86546 3502 86548 3554
rect 86492 3490 86548 3502
rect 86156 3332 86212 3342
rect 86156 3238 86212 3276
rect 87500 800 87556 3612
rect 88172 3554 88228 4398
rect 88284 4452 88340 4844
rect 88284 4386 88340 4396
rect 89068 4898 89124 4910
rect 89068 4846 89070 4898
rect 89122 4846 89124 4898
rect 89068 3780 89124 4846
rect 89292 4452 89348 4462
rect 89292 4358 89348 4396
rect 89628 4450 89684 4462
rect 89628 4398 89630 4450
rect 89682 4398 89684 4450
rect 89068 3714 89124 3724
rect 88732 3668 88788 3678
rect 88732 3574 88788 3612
rect 89180 3668 89236 3678
rect 88172 3502 88174 3554
rect 88226 3502 88228 3554
rect 88172 3490 88228 3502
rect 89180 800 89236 3612
rect 89628 3556 89684 4398
rect 90188 4450 90244 5180
rect 90188 4398 90190 4450
rect 90242 4398 90244 4450
rect 90188 4386 90244 4398
rect 90300 5234 90356 8876
rect 90300 5182 90302 5234
rect 90354 5182 90356 5234
rect 90300 4452 90356 5182
rect 90748 5236 90804 9884
rect 93262 8652 93526 8662
rect 93318 8596 93366 8652
rect 93422 8596 93470 8652
rect 93262 8586 93526 8596
rect 90748 5104 90804 5180
rect 91532 7252 91588 7262
rect 91532 4788 91588 7196
rect 93262 7084 93526 7094
rect 93318 7028 93366 7084
rect 93422 7028 93470 7084
rect 93262 7018 93526 7028
rect 97356 6020 97412 6030
rect 96460 5794 96516 5806
rect 96460 5742 96462 5794
rect 96514 5742 96516 5794
rect 96460 5684 96516 5742
rect 96460 5618 96516 5628
rect 93262 5516 93526 5526
rect 93318 5460 93366 5516
rect 93422 5460 93470 5516
rect 93262 5450 93526 5460
rect 96460 5460 96516 5470
rect 96236 5348 96292 5358
rect 96236 5254 96292 5292
rect 91532 4722 91588 4732
rect 94108 5236 94164 5246
rect 90300 4386 90356 4396
rect 90524 4452 90580 4462
rect 90524 4358 90580 4396
rect 91084 4452 91140 4462
rect 91084 4338 91140 4396
rect 93996 4452 94052 4462
rect 93996 4358 94052 4396
rect 91084 4286 91086 4338
rect 91138 4286 91140 4338
rect 91084 4274 91140 4286
rect 90860 4228 90916 4238
rect 90524 3668 90580 3678
rect 90524 3574 90580 3612
rect 89852 3556 89908 3566
rect 89628 3554 89908 3556
rect 89628 3502 89854 3554
rect 89906 3502 89908 3554
rect 89628 3500 89908 3502
rect 89852 3490 89908 3500
rect 90860 800 90916 4172
rect 91756 4228 91812 4238
rect 91756 4134 91812 4172
rect 93262 3948 93526 3958
rect 93318 3892 93366 3948
rect 93422 3892 93470 3948
rect 93262 3882 93526 3892
rect 94108 3666 94164 5180
rect 95452 5124 95508 5134
rect 95452 5030 95508 5068
rect 95900 5122 95956 5134
rect 95900 5070 95902 5122
rect 95954 5070 95956 5122
rect 95116 5012 95172 5022
rect 94668 5010 95172 5012
rect 94668 4958 95118 5010
rect 95170 4958 95172 5010
rect 94668 4956 95172 4958
rect 94556 4900 94612 4910
rect 94668 4900 94724 4956
rect 95116 4946 95172 4956
rect 94556 4898 94724 4900
rect 94556 4846 94558 4898
rect 94610 4846 94724 4898
rect 94556 4844 94724 4846
rect 94556 4834 94612 4844
rect 94108 3614 94110 3666
rect 94162 3614 94164 3666
rect 94108 3602 94164 3614
rect 94220 4452 94276 4462
rect 92316 3444 92372 3454
rect 92876 3444 92932 3454
rect 92316 3442 92932 3444
rect 92316 3390 92318 3442
rect 92370 3390 92878 3442
rect 92930 3390 92932 3442
rect 92316 3388 92932 3390
rect 92316 3378 92372 3388
rect 92540 800 92596 3388
rect 92876 3378 92932 3388
rect 94220 800 94276 4396
rect 94556 4452 94612 4462
rect 94556 4358 94612 4396
rect 94668 1652 94724 4844
rect 95900 4226 95956 5070
rect 96460 4562 96516 5404
rect 97020 5460 97076 5470
rect 97020 5010 97076 5404
rect 97020 4958 97022 5010
rect 97074 4958 97076 5010
rect 97020 4946 97076 4958
rect 97132 5124 97188 5134
rect 97356 5124 97412 5964
rect 97468 6018 97524 6030
rect 97468 5966 97470 6018
rect 97522 5966 97524 6018
rect 97468 5684 97524 5966
rect 97916 6020 97972 6030
rect 97916 5926 97972 5964
rect 97468 5618 97524 5628
rect 98028 5348 98084 11116
rect 98476 6130 98532 12124
rect 98476 6078 98478 6130
rect 98530 6078 98532 6130
rect 98476 6066 98532 6078
rect 99036 6020 99092 6030
rect 99036 5794 99092 5964
rect 99036 5742 99038 5794
rect 99090 5742 99092 5794
rect 98140 5684 98196 5694
rect 98140 5682 98308 5684
rect 98140 5630 98142 5682
rect 98194 5630 98308 5682
rect 98140 5628 98308 5630
rect 98140 5618 98196 5628
rect 98140 5348 98196 5358
rect 98028 5346 98196 5348
rect 98028 5294 98142 5346
rect 98194 5294 98196 5346
rect 98028 5292 98196 5294
rect 98140 5282 98196 5292
rect 97188 5122 97412 5124
rect 97188 5070 97358 5122
rect 97410 5070 97412 5122
rect 97188 5068 97412 5070
rect 96460 4510 96462 4562
rect 96514 4510 96516 4562
rect 96460 4498 96516 4510
rect 97132 4562 97188 5068
rect 97356 5058 97412 5068
rect 97804 5122 97860 5134
rect 97804 5070 97806 5122
rect 97858 5070 97860 5122
rect 97132 4510 97134 4562
rect 97186 4510 97188 4562
rect 97132 4498 97188 4510
rect 95900 4174 95902 4226
rect 95954 4174 95956 4226
rect 95900 4162 95956 4174
rect 97580 3668 97636 3678
rect 97804 3668 97860 5070
rect 97580 3666 97860 3668
rect 97580 3614 97582 3666
rect 97634 3614 97860 3666
rect 97580 3612 97860 3614
rect 98028 4450 98084 4462
rect 98028 4398 98030 4450
rect 98082 4398 98084 4450
rect 97580 3602 97636 3612
rect 95228 3444 95284 3482
rect 95228 3378 95284 3388
rect 95900 3444 95956 3454
rect 94668 1586 94724 1596
rect 95900 800 95956 3388
rect 96236 3444 96292 3482
rect 96236 3378 96292 3388
rect 97580 3444 97636 3454
rect 97580 800 97636 3388
rect 98028 3444 98084 4398
rect 98252 4228 98308 5628
rect 99036 5124 99092 5742
rect 99484 5794 99540 5806
rect 99484 5742 99486 5794
rect 99538 5742 99540 5794
rect 99260 5124 99316 5134
rect 99036 5068 99260 5124
rect 99260 5030 99316 5068
rect 99484 5124 99540 5742
rect 100044 5346 100100 12796
rect 100492 12402 100548 14252
rect 101164 12852 101220 12862
rect 101164 12758 101220 12796
rect 101500 12852 101556 12862
rect 101500 12758 101556 12796
rect 100492 12350 100494 12402
rect 100546 12350 100548 12402
rect 100492 12338 100548 12350
rect 100156 12180 100212 12190
rect 100156 12086 100212 12124
rect 101164 11282 101220 11294
rect 101164 11230 101166 11282
rect 101218 11230 101220 11282
rect 100492 11172 100548 11182
rect 100492 11078 100548 11116
rect 101164 11172 101220 11230
rect 101164 11106 101220 11116
rect 101500 11172 101556 11182
rect 101500 11078 101556 11116
rect 101948 10612 102004 10622
rect 101500 7700 101556 7710
rect 100044 5294 100046 5346
rect 100098 5294 100100 5346
rect 100044 5282 100100 5294
rect 101164 6578 101220 6590
rect 101164 6526 101166 6578
rect 101218 6526 101220 6578
rect 101164 5348 101220 6526
rect 101500 6578 101556 7644
rect 101500 6526 101502 6578
rect 101554 6526 101556 6578
rect 101500 6514 101556 6526
rect 101948 6130 102004 10556
rect 103292 6580 103348 6590
rect 101948 6078 101950 6130
rect 102002 6078 102004 6130
rect 101948 6020 102004 6078
rect 102956 6578 103348 6580
rect 102956 6526 103294 6578
rect 103346 6526 103348 6578
rect 102956 6524 103348 6526
rect 101948 5954 102004 5964
rect 102732 6020 102788 6030
rect 102732 5926 102788 5964
rect 101164 5282 101220 5292
rect 101388 5908 101444 5918
rect 99484 5058 99540 5068
rect 99708 5124 99764 5134
rect 101052 5124 101108 5134
rect 99708 5122 99876 5124
rect 99708 5070 99710 5122
rect 99762 5070 99876 5122
rect 99708 5068 99876 5070
rect 99708 5058 99764 5068
rect 98252 4162 98308 4172
rect 98588 5012 98644 5022
rect 98588 3666 98644 4956
rect 98924 5012 98980 5022
rect 98924 4918 98980 4956
rect 99036 4228 99092 4238
rect 99036 4134 99092 4172
rect 98588 3614 98590 3666
rect 98642 3614 98644 3666
rect 98588 3602 98644 3614
rect 99820 3666 99876 5068
rect 101052 5030 101108 5068
rect 101276 4452 101332 4462
rect 100940 4450 101332 4452
rect 100940 4398 101278 4450
rect 101330 4398 101332 4450
rect 100940 4396 101332 4398
rect 100716 4228 100772 4238
rect 100940 4228 100996 4396
rect 101276 4386 101332 4396
rect 100716 4226 100996 4228
rect 100716 4174 100718 4226
rect 100770 4174 100996 4226
rect 100716 4172 100996 4174
rect 100716 4162 100772 4172
rect 99820 3614 99822 3666
rect 99874 3614 99876 3666
rect 99820 3602 99876 3614
rect 98028 3350 98084 3388
rect 99148 3444 99204 3454
rect 99260 3444 99316 3454
rect 99148 3442 99260 3444
rect 99148 3390 99150 3442
rect 99202 3390 99260 3442
rect 99148 3388 99260 3390
rect 99148 3378 99204 3388
rect 99260 800 99316 3388
rect 100828 3444 100884 3454
rect 100828 3350 100884 3388
rect 100940 800 100996 4172
rect 101388 3780 101444 5852
rect 102172 5908 102228 5918
rect 101500 5794 101556 5806
rect 101500 5742 101502 5794
rect 101554 5742 101556 5794
rect 101500 5012 101556 5742
rect 102172 5122 102228 5852
rect 102620 5908 102676 5918
rect 102620 5814 102676 5852
rect 102956 5346 103012 6524
rect 103292 6514 103348 6524
rect 103628 6578 103684 15820
rect 104188 6580 104244 6590
rect 103628 6526 103630 6578
rect 103682 6526 103684 6578
rect 103628 6514 103684 6526
rect 103740 6578 104244 6580
rect 103740 6526 104190 6578
rect 104242 6526 104244 6578
rect 103740 6524 104244 6526
rect 103740 6130 103796 6524
rect 104188 6514 104244 6524
rect 104524 6578 104580 16828
rect 105868 10836 105924 10846
rect 105868 8428 105924 10780
rect 105532 8372 105924 8428
rect 105532 7698 105588 8372
rect 105532 7646 105534 7698
rect 105586 7646 105588 7698
rect 105532 7634 105588 7646
rect 105308 7474 105364 7486
rect 105308 7422 105310 7474
rect 105362 7422 105364 7474
rect 105196 6580 105252 6590
rect 104524 6526 104526 6578
rect 104578 6526 104580 6578
rect 104524 6514 104580 6526
rect 104860 6578 105252 6580
rect 104860 6526 105198 6578
rect 105250 6526 105252 6578
rect 104860 6524 105252 6526
rect 103740 6078 103742 6130
rect 103794 6078 103796 6130
rect 103740 6066 103796 6078
rect 103740 5908 103796 5918
rect 102956 5294 102958 5346
rect 103010 5294 103012 5346
rect 102956 5282 103012 5294
rect 103404 5682 103460 5694
rect 103404 5630 103406 5682
rect 103458 5630 103460 5682
rect 102172 5070 102174 5122
rect 102226 5070 102228 5122
rect 102172 5058 102228 5070
rect 102620 5122 102676 5134
rect 102620 5070 102622 5122
rect 102674 5070 102676 5122
rect 101836 5012 101892 5022
rect 101500 5010 101892 5012
rect 101500 4958 101838 5010
rect 101890 4958 101892 5010
rect 101500 4956 101892 4958
rect 101388 3714 101444 3724
rect 101836 2324 101892 4956
rect 102620 4226 102676 5070
rect 102620 4174 102622 4226
rect 102674 4174 102676 4226
rect 102620 4162 102676 4174
rect 103292 4226 103348 4238
rect 103292 4174 103294 4226
rect 103346 4174 103348 4226
rect 103292 4004 103348 4174
rect 103292 3938 103348 3948
rect 103404 3668 103460 5630
rect 103740 5348 103796 5852
rect 103740 5122 103796 5292
rect 104412 5794 104468 5806
rect 104412 5742 104414 5794
rect 104466 5742 104468 5794
rect 103740 5070 103742 5122
rect 103794 5070 103796 5122
rect 103740 5058 103796 5070
rect 103852 5124 103908 5134
rect 103852 4226 103908 5068
rect 103964 5012 104020 5022
rect 103964 4918 104020 4956
rect 104412 5012 104468 5742
rect 104860 5346 104916 6524
rect 105196 6514 105252 6524
rect 105308 6130 105364 7422
rect 105532 7364 105588 7374
rect 105532 6578 105588 7308
rect 106652 7364 106708 17388
rect 106652 7298 106708 7308
rect 107772 15092 107828 15102
rect 105532 6526 105534 6578
rect 105586 6526 105588 6578
rect 105532 6514 105588 6526
rect 105308 6078 105310 6130
rect 105362 6078 105364 6130
rect 105308 6066 105364 6078
rect 105980 6466 106036 6478
rect 105980 6414 105982 6466
rect 106034 6414 106036 6466
rect 104860 5294 104862 5346
rect 104914 5294 104916 5346
rect 104860 5282 104916 5294
rect 105644 5684 105700 5694
rect 105980 5684 106036 6414
rect 106988 6132 107044 6142
rect 106204 6130 107044 6132
rect 106204 6078 106990 6130
rect 107042 6078 107044 6130
rect 106204 6076 107044 6078
rect 106204 6020 106260 6076
rect 106988 6066 107044 6076
rect 105644 5682 106036 5684
rect 105644 5630 105646 5682
rect 105698 5630 106036 5682
rect 105644 5628 106036 5630
rect 106092 6018 106260 6020
rect 106092 5966 106206 6018
rect 106258 5966 106260 6018
rect 106092 5964 106260 5966
rect 105644 5236 105700 5628
rect 105644 5170 105700 5180
rect 105868 5348 105924 5358
rect 104412 4946 104468 4956
rect 104524 5122 104580 5134
rect 104524 5070 104526 5122
rect 104578 5070 104580 5122
rect 103852 4174 103854 4226
rect 103906 4174 103908 4226
rect 103852 4162 103908 4174
rect 104300 4338 104356 4350
rect 104300 4286 104302 4338
rect 104354 4286 104356 4338
rect 104300 4004 104356 4286
rect 104524 4228 104580 5070
rect 105868 5122 105924 5292
rect 105868 5070 105870 5122
rect 105922 5070 105924 5122
rect 105644 5010 105700 5022
rect 105644 4958 105646 5010
rect 105698 4958 105700 5010
rect 105644 4788 105700 4958
rect 105644 4722 105700 4732
rect 105196 4228 105252 4238
rect 104524 4226 105252 4228
rect 104524 4174 105198 4226
rect 105250 4174 105252 4226
rect 104524 4172 105252 4174
rect 105196 4162 105252 4172
rect 104300 3938 104356 3948
rect 103740 3668 103796 3678
rect 103404 3666 103796 3668
rect 103404 3614 103742 3666
rect 103794 3614 103796 3666
rect 103404 3612 103796 3614
rect 103740 3602 103796 3612
rect 105868 3666 105924 5070
rect 105868 3614 105870 3666
rect 105922 3614 105924 3666
rect 105868 3602 105924 3614
rect 104300 3556 104356 3566
rect 101836 2258 101892 2268
rect 103068 3444 103124 3454
rect 103068 2212 103124 3388
rect 102620 2156 103124 2212
rect 102620 800 102676 2156
rect 104300 800 104356 3500
rect 104748 3444 104804 3454
rect 104748 3350 104804 3388
rect 105980 3444 106036 3454
rect 105980 800 106036 3388
rect 106092 2436 106148 5964
rect 106204 5954 106260 5964
rect 106428 5906 106484 5918
rect 106428 5854 106430 5906
rect 106482 5854 106484 5906
rect 106428 5684 106484 5854
rect 107436 5794 107492 5806
rect 107436 5742 107438 5794
rect 107490 5742 107492 5794
rect 106764 5684 106820 5694
rect 106428 5682 106820 5684
rect 106428 5630 106766 5682
rect 106818 5630 106820 5682
rect 106428 5628 106820 5630
rect 106764 5618 106820 5628
rect 107436 5682 107492 5742
rect 107436 5630 107438 5682
rect 107490 5630 107492 5682
rect 107436 5236 107492 5630
rect 107436 5180 107604 5236
rect 106428 5122 106484 5134
rect 106428 5070 106430 5122
rect 106482 5070 106484 5122
rect 106204 4450 106260 4462
rect 106204 4398 106206 4450
rect 106258 4398 106260 4450
rect 106204 3556 106260 4398
rect 106204 3490 106260 3500
rect 106316 4004 106372 4014
rect 106316 3554 106372 3948
rect 106428 3668 106484 5070
rect 106764 5012 106820 5022
rect 107436 5012 107492 5022
rect 106764 5010 107492 5012
rect 106764 4958 106766 5010
rect 106818 4958 107438 5010
rect 107490 4958 107492 5010
rect 106764 4956 107492 4958
rect 106764 4946 106820 4956
rect 107436 4946 107492 4956
rect 107100 4788 107156 4798
rect 107548 4788 107604 5180
rect 107772 5010 107828 15036
rect 109116 6804 109172 6814
rect 109116 6244 109172 6748
rect 110460 6690 110516 6702
rect 110460 6638 110462 6690
rect 110514 6638 110516 6690
rect 109116 6130 109172 6188
rect 109116 6078 109118 6130
rect 109170 6078 109172 6130
rect 109116 6066 109172 6078
rect 109900 6244 109956 6254
rect 109900 6018 109956 6188
rect 109900 5966 109902 6018
rect 109954 5966 109956 6018
rect 109900 5954 109956 5966
rect 109788 5908 109844 5918
rect 107772 4958 107774 5010
rect 107826 4958 107828 5010
rect 107772 4946 107828 4958
rect 107884 5794 107940 5806
rect 107884 5742 107886 5794
rect 107938 5742 107940 5794
rect 107100 4562 107156 4732
rect 107100 4510 107102 4562
rect 107154 4510 107156 4562
rect 107100 4498 107156 4510
rect 107436 4732 107604 4788
rect 107436 3892 107492 4732
rect 107436 3826 107492 3836
rect 106428 3602 106484 3612
rect 107660 3668 107716 3678
rect 107660 3574 107716 3612
rect 106316 3502 106318 3554
rect 106370 3502 106372 3554
rect 106316 3490 106372 3502
rect 106764 3556 106820 3566
rect 106764 3462 106820 3500
rect 107884 3444 107940 5742
rect 108780 5796 108836 5806
rect 108780 5794 109284 5796
rect 108780 5742 108782 5794
rect 108834 5742 109284 5794
rect 108780 5740 109284 5742
rect 108780 5730 108836 5740
rect 109228 5010 109284 5740
rect 109564 5124 109620 5134
rect 109564 5030 109620 5068
rect 109788 5124 109844 5852
rect 110460 5908 110516 6638
rect 110908 6130 110964 18172
rect 111672 17276 111936 17286
rect 111728 17220 111776 17276
rect 111832 17220 111880 17276
rect 111672 17210 111936 17220
rect 111672 15708 111936 15718
rect 111728 15652 111776 15708
rect 111832 15652 111880 15708
rect 111672 15642 111936 15652
rect 111672 14140 111936 14150
rect 111728 14084 111776 14140
rect 111832 14084 111880 14140
rect 111672 14074 111936 14084
rect 111672 12572 111936 12582
rect 111728 12516 111776 12572
rect 111832 12516 111880 12572
rect 111672 12506 111936 12516
rect 111672 11004 111936 11014
rect 111728 10948 111776 11004
rect 111832 10948 111880 11004
rect 111672 10938 111936 10948
rect 111672 9436 111936 9446
rect 111728 9380 111776 9436
rect 111832 9380 111880 9436
rect 111672 9370 111936 9380
rect 111672 7868 111936 7878
rect 111728 7812 111776 7868
rect 111832 7812 111880 7868
rect 111672 7802 111936 7812
rect 110908 6078 110910 6130
rect 110962 6078 110964 6130
rect 110908 6066 110964 6078
rect 111020 6468 111076 6478
rect 111468 6468 111524 6478
rect 111020 6466 111524 6468
rect 111020 6414 111022 6466
rect 111074 6414 111470 6466
rect 111522 6414 111524 6466
rect 111020 6412 111524 6414
rect 110460 5842 110516 5852
rect 110572 5684 110628 5694
rect 110124 5682 110628 5684
rect 110124 5630 110574 5682
rect 110626 5630 110628 5682
rect 110124 5628 110628 5630
rect 109788 5058 109844 5068
rect 110012 5122 110068 5134
rect 110012 5070 110014 5122
rect 110066 5070 110068 5122
rect 109228 4958 109230 5010
rect 109282 4958 109284 5010
rect 108220 4898 108276 4910
rect 108220 4846 108222 4898
rect 108274 4846 108276 4898
rect 107884 3378 107940 3388
rect 107996 4452 108052 4462
rect 108220 4452 108276 4846
rect 107996 4450 108276 4452
rect 107996 4398 107998 4450
rect 108050 4398 108276 4450
rect 107996 4396 108276 4398
rect 108332 4900 108388 4910
rect 107996 3108 108052 4396
rect 106092 2370 106148 2380
rect 107660 3052 108052 3108
rect 107660 800 107716 3052
rect 108332 2548 108388 4844
rect 109228 4564 109284 4958
rect 109228 4498 109284 4508
rect 109340 4228 109396 4238
rect 110012 4228 110068 5070
rect 109340 4226 110068 4228
rect 109340 4174 109342 4226
rect 109394 4174 110068 4226
rect 109340 4172 110068 4174
rect 110124 4226 110180 5628
rect 110572 5618 110628 5628
rect 110124 4174 110126 4226
rect 110178 4174 110180 4226
rect 109340 4162 109396 4172
rect 110124 4162 110180 4174
rect 110348 4898 110404 4910
rect 110348 4846 110350 4898
rect 110402 4846 110404 4898
rect 109564 4004 109620 4014
rect 109340 3668 109396 3678
rect 108668 3444 108724 3454
rect 108668 3350 108724 3388
rect 108332 2482 108388 2492
rect 109340 800 109396 3612
rect 109564 3666 109620 3948
rect 109564 3614 109566 3666
rect 109618 3614 109620 3666
rect 109564 3602 109620 3614
rect 110348 3554 110404 4846
rect 110908 4450 110964 4462
rect 110908 4398 110910 4450
rect 110962 4398 110964 4450
rect 110908 4228 110964 4398
rect 110908 3668 110964 4172
rect 111020 4004 111076 6412
rect 111468 6402 111524 6412
rect 112700 6466 112756 6478
rect 112700 6414 112702 6466
rect 112754 6414 112756 6466
rect 111672 6300 111936 6310
rect 111728 6244 111776 6300
rect 111832 6244 111880 6300
rect 111672 6234 111936 6244
rect 112028 6018 112084 6030
rect 112028 5966 112030 6018
rect 112082 5966 112084 6018
rect 111804 5906 111860 5918
rect 111804 5854 111806 5906
rect 111858 5854 111860 5906
rect 111804 5348 111860 5854
rect 112028 5796 112084 5966
rect 112028 5730 112084 5740
rect 112252 5348 112308 5358
rect 111804 5346 112308 5348
rect 111804 5294 112254 5346
rect 112306 5294 112308 5346
rect 111804 5292 112308 5294
rect 112252 5282 112308 5292
rect 111468 5124 111524 5134
rect 111468 5030 111524 5068
rect 111916 5124 111972 5134
rect 111916 5122 112084 5124
rect 111916 5070 111918 5122
rect 111970 5070 112084 5122
rect 111916 5068 112084 5070
rect 111916 5058 111972 5068
rect 111020 3938 111076 3948
rect 111132 5010 111188 5022
rect 111132 4958 111134 5010
rect 111186 4958 111188 5010
rect 110908 3602 110964 3612
rect 110348 3502 110350 3554
rect 110402 3502 110404 3554
rect 110348 3490 110404 3502
rect 111020 3556 111076 3566
rect 110684 3330 110740 3342
rect 110684 3278 110686 3330
rect 110738 3278 110740 3330
rect 110684 2548 110740 3278
rect 110684 2482 110740 2492
rect 111020 800 111076 3500
rect 111132 2884 111188 4958
rect 111672 4732 111936 4742
rect 111728 4676 111776 4732
rect 111832 4676 111880 4732
rect 111672 4666 111936 4676
rect 111804 4228 111860 4238
rect 111804 4134 111860 4172
rect 111804 3668 111860 3678
rect 112028 3668 112084 5068
rect 112700 5012 112756 6414
rect 113484 6130 113540 22092
rect 114268 20580 114324 20590
rect 114268 18676 114324 20524
rect 114268 18610 114324 18620
rect 115836 18340 115892 18350
rect 115836 15092 115892 18284
rect 115836 15026 115892 15036
rect 117404 14420 117460 14430
rect 113484 6078 113486 6130
rect 113538 6078 113540 6130
rect 113484 6066 113540 6078
rect 115276 9156 115332 9166
rect 115276 6130 115332 9100
rect 117068 6580 117124 6590
rect 115276 6078 115278 6130
rect 115330 6078 115332 6130
rect 115276 6020 115332 6078
rect 116172 6578 117124 6580
rect 116172 6526 117070 6578
rect 117122 6526 117124 6578
rect 116172 6524 117124 6526
rect 115276 5954 115332 5964
rect 116060 6020 116116 6030
rect 116060 5926 116116 5964
rect 113260 5908 113316 5918
rect 115388 5908 115444 5918
rect 113260 5906 114212 5908
rect 113260 5854 113262 5906
rect 113314 5854 114212 5906
rect 113260 5852 114212 5854
rect 113260 5842 113316 5852
rect 114156 5346 114212 5852
rect 114156 5294 114158 5346
rect 114210 5294 114212 5346
rect 114156 5282 114212 5294
rect 114716 5794 114772 5806
rect 114716 5742 114718 5794
rect 114770 5742 114772 5794
rect 113148 5124 113204 5134
rect 113148 5030 113204 5068
rect 113820 5122 113876 5134
rect 113820 5070 113822 5122
rect 113874 5070 113876 5122
rect 113036 5012 113092 5022
rect 112700 5010 113092 5012
rect 112700 4958 113038 5010
rect 113090 4958 113092 5010
rect 112700 4956 113092 4958
rect 111804 3666 112084 3668
rect 111804 3614 111806 3666
rect 111858 3614 112084 3666
rect 111804 3612 112084 3614
rect 112252 4226 112308 4238
rect 112252 4174 112254 4226
rect 112306 4174 112308 4226
rect 111804 3602 111860 3612
rect 111672 3164 111936 3174
rect 111728 3108 111776 3164
rect 111832 3108 111880 3164
rect 111672 3098 111936 3108
rect 111132 2818 111188 2828
rect 112252 2884 112308 4174
rect 112588 3556 112644 3566
rect 112588 3442 112644 3500
rect 112588 3390 112590 3442
rect 112642 3390 112644 3442
rect 112588 3378 112644 3390
rect 112700 3444 112756 3454
rect 112252 2818 112308 2828
rect 112700 800 112756 3388
rect 113036 1092 113092 4956
rect 113260 4450 113316 4462
rect 113260 4398 113262 4450
rect 113314 4398 113316 4450
rect 113260 3444 113316 4398
rect 113820 4228 113876 5070
rect 114716 5012 114772 5742
rect 115388 5122 115444 5852
rect 116172 5346 116228 6524
rect 117068 6514 117124 6524
rect 117404 6578 117460 14364
rect 117964 7588 118020 7598
rect 117964 6692 118020 7532
rect 119196 6804 119252 24556
rect 119196 6738 119252 6748
rect 119308 7028 119364 7038
rect 117964 6690 118132 6692
rect 117964 6638 117966 6690
rect 118018 6638 118132 6690
rect 117964 6636 118132 6638
rect 117964 6626 118020 6636
rect 117404 6526 117406 6578
rect 117458 6526 117460 6578
rect 117404 6514 117460 6526
rect 116508 6020 116564 6030
rect 116508 5926 116564 5964
rect 117740 6020 117796 6030
rect 117740 5908 117796 5964
rect 118076 6018 118132 6636
rect 118076 5966 118078 6018
rect 118130 5966 118132 6018
rect 118076 5954 118132 5966
rect 117964 5908 118020 5918
rect 117740 5906 118020 5908
rect 117740 5854 117966 5906
rect 118018 5854 118020 5906
rect 117740 5852 118020 5854
rect 116172 5294 116174 5346
rect 116226 5294 116228 5346
rect 116172 5282 116228 5294
rect 116732 5682 116788 5694
rect 116732 5630 116734 5682
rect 116786 5630 116788 5682
rect 115388 5070 115390 5122
rect 115442 5070 115444 5122
rect 115388 5058 115444 5070
rect 115836 5122 115892 5134
rect 115836 5070 115838 5122
rect 115890 5070 115892 5122
rect 115052 5012 115108 5022
rect 114716 5010 115108 5012
rect 114716 4958 115054 5010
rect 115106 4958 115108 5010
rect 114716 4956 115108 4958
rect 113820 4162 113876 4172
rect 114380 4228 114436 4238
rect 114380 4134 114436 4172
rect 113484 3556 113540 3566
rect 113484 3462 113540 3500
rect 113260 3378 113316 3388
rect 113932 3444 113988 3454
rect 113932 3350 113988 3388
rect 114828 3444 114884 3454
rect 114828 2212 114884 3388
rect 113036 1026 113092 1036
rect 114380 2156 114884 2212
rect 114380 800 114436 2156
rect 115052 1540 115108 4956
rect 115724 5012 115780 5022
rect 115388 4228 115444 4238
rect 115388 4134 115444 4172
rect 115724 4226 115780 4956
rect 115724 4174 115726 4226
rect 115778 4174 115780 4226
rect 115612 3444 115668 3454
rect 115612 3350 115668 3388
rect 115724 2772 115780 4174
rect 115836 3668 115892 5070
rect 116396 4452 116452 4462
rect 115836 3602 115892 3612
rect 116060 4450 116452 4452
rect 116060 4398 116398 4450
rect 116450 4398 116452 4450
rect 116060 4396 116452 4398
rect 116060 4228 116116 4396
rect 116396 4386 116452 4396
rect 115724 2706 115780 2716
rect 115052 1474 115108 1484
rect 116060 800 116116 4172
rect 116732 4228 116788 5630
rect 117068 5682 117124 5694
rect 117068 5630 117070 5682
rect 117122 5630 117124 5682
rect 117068 4900 117124 5630
rect 117180 5012 117236 5022
rect 117180 4918 117236 4956
rect 117740 5010 117796 5852
rect 117964 5842 118020 5852
rect 119084 5908 119140 5918
rect 119084 5814 119140 5852
rect 118748 5682 118804 5694
rect 118748 5630 118750 5682
rect 118802 5630 118804 5682
rect 117740 4958 117742 5010
rect 117794 4958 117796 5010
rect 117068 4834 117124 4844
rect 116732 4162 116788 4172
rect 117516 4228 117572 4238
rect 117516 4134 117572 4172
rect 116732 3668 116788 3678
rect 116732 3574 116788 3612
rect 117628 3668 117684 3678
rect 117740 3668 117796 4958
rect 117964 5122 118020 5134
rect 117964 5070 117966 5122
rect 118018 5070 118020 5122
rect 117964 4228 118020 5070
rect 118300 5012 118356 5022
rect 118300 4918 118356 4956
rect 118300 4228 118356 4238
rect 117964 4226 118356 4228
rect 117964 4174 118302 4226
rect 118354 4174 118356 4226
rect 117964 4172 118356 4174
rect 118300 4162 118356 4172
rect 117628 3666 117796 3668
rect 117628 3614 117630 3666
rect 117682 3614 117796 3666
rect 117628 3612 117796 3614
rect 118076 3892 118132 3902
rect 117628 3602 117684 3612
rect 118076 3554 118132 3836
rect 118748 3668 118804 5630
rect 118972 5010 119028 5022
rect 118972 4958 118974 5010
rect 119026 4958 119028 5010
rect 118972 4900 119028 4958
rect 119308 5010 119364 6972
rect 120092 6130 120148 25116
rect 121772 23716 121828 23726
rect 121772 7028 121828 23660
rect 121772 6962 121828 6972
rect 122108 10724 122164 10734
rect 120092 6078 120094 6130
rect 120146 6078 120148 6130
rect 120092 6066 120148 6078
rect 120204 6804 120260 6814
rect 119756 5908 119812 5918
rect 119756 5814 119812 5852
rect 119308 4958 119310 5010
rect 119362 4958 119364 5010
rect 119308 4946 119364 4958
rect 119868 5012 119924 5022
rect 119868 4918 119924 4956
rect 120204 5010 120260 6748
rect 122108 6130 122164 10668
rect 122108 6078 122110 6130
rect 122162 6078 122164 6130
rect 122108 6020 122164 6078
rect 122668 7812 122724 7822
rect 122668 6132 122724 7756
rect 122668 6066 122724 6076
rect 122108 5954 122164 5964
rect 122892 6020 122948 6030
rect 122892 5926 122948 5964
rect 123340 6018 123396 6030
rect 123340 5966 123342 6018
rect 123394 5966 123396 6018
rect 123340 5796 123396 5966
rect 123900 5908 123956 5918
rect 123900 5814 123956 5852
rect 123396 5740 123508 5796
rect 123340 5730 123396 5740
rect 122332 5236 122388 5246
rect 122332 5122 122388 5180
rect 123452 5236 123508 5740
rect 122332 5070 122334 5122
rect 122386 5070 122388 5122
rect 122332 5058 122388 5070
rect 122780 5122 122836 5134
rect 122780 5070 122782 5122
rect 122834 5070 122836 5122
rect 121996 5012 122052 5022
rect 120204 4958 120206 5010
rect 120258 4958 120260 5010
rect 120204 4946 120260 4958
rect 121436 5010 122052 5012
rect 121436 4958 121998 5010
rect 122050 4958 122052 5010
rect 121436 4956 122052 4958
rect 121436 4900 121492 4956
rect 121996 4946 122052 4956
rect 118972 4834 119028 4844
rect 121324 4898 121492 4900
rect 121324 4846 121438 4898
rect 121490 4846 121492 4898
rect 121324 4844 121492 4846
rect 120204 4564 120260 4574
rect 119308 4452 119364 4462
rect 118748 3602 118804 3612
rect 119196 4450 119364 4452
rect 119196 4398 119310 4450
rect 119362 4398 119364 4450
rect 119196 4396 119364 4398
rect 118076 3502 118078 3554
rect 118130 3502 118132 3554
rect 118076 3490 118132 3502
rect 117740 3444 117796 3454
rect 117740 800 117796 3388
rect 118524 3444 118580 3454
rect 118524 3350 118580 3388
rect 119196 3444 119252 4396
rect 119308 4386 119364 4396
rect 120204 3892 120260 4508
rect 120204 3826 120260 3836
rect 119644 3668 119700 3678
rect 119644 3574 119700 3612
rect 120652 3668 120708 3678
rect 119196 3378 119252 3388
rect 119420 3444 119476 3454
rect 119420 800 119476 3388
rect 120652 3444 120708 3612
rect 120652 3350 120708 3388
rect 121100 3444 121156 3454
rect 121100 800 121156 3388
rect 121324 1316 121380 4844
rect 121436 4834 121492 4844
rect 121436 4450 121492 4462
rect 121436 4398 121438 4450
rect 121490 4398 121492 4450
rect 121436 3444 121492 4398
rect 122780 4226 122836 5070
rect 123116 5012 123172 5022
rect 123116 4918 123172 4956
rect 123452 4562 123508 5180
rect 123452 4510 123454 4562
rect 123506 4510 123508 4562
rect 123452 4498 123508 4510
rect 123564 5682 123620 5694
rect 123564 5630 123566 5682
rect 123618 5630 123620 5682
rect 122780 4174 122782 4226
rect 122834 4174 122836 4226
rect 122780 4162 122836 4174
rect 121548 3668 121604 3678
rect 121548 3574 121604 3612
rect 123564 3666 123620 5630
rect 123788 5012 123844 5022
rect 123788 4918 123844 4956
rect 124124 5010 124180 26908
rect 124348 6466 124404 6478
rect 124348 6414 124350 6466
rect 124402 6414 124404 6466
rect 124348 5796 124404 6414
rect 124908 6130 124964 27692
rect 124908 6078 124910 6130
rect 124962 6078 124964 6130
rect 124908 6066 124964 6078
rect 126028 22932 126084 22942
rect 126028 6130 126084 22876
rect 126028 6078 126030 6130
rect 126082 6078 126084 6130
rect 126028 6066 126084 6078
rect 126924 8484 126980 8494
rect 124572 5908 124628 5918
rect 124572 5814 124628 5852
rect 125804 5908 125860 5918
rect 125804 5906 126308 5908
rect 125804 5854 125806 5906
rect 125858 5854 126308 5906
rect 125804 5852 126308 5854
rect 125804 5842 125860 5852
rect 124348 5730 124404 5740
rect 125468 5796 125524 5806
rect 125468 5122 125524 5740
rect 126252 5346 126308 5852
rect 126252 5294 126254 5346
rect 126306 5294 126308 5346
rect 126252 5282 126308 5294
rect 126588 5796 126644 5806
rect 125468 5070 125470 5122
rect 125522 5070 125524 5122
rect 125468 5058 125524 5070
rect 125916 5122 125972 5134
rect 125916 5070 125918 5122
rect 125970 5070 125972 5122
rect 124124 4958 124126 5010
rect 124178 4958 124180 5010
rect 124124 4946 124180 4958
rect 124908 5012 124964 5022
rect 124796 4452 124852 4462
rect 124460 4450 124852 4452
rect 124460 4398 124798 4450
rect 124850 4398 124852 4450
rect 124460 4396 124852 4398
rect 124236 4228 124292 4238
rect 124460 4228 124516 4396
rect 124796 4386 124852 4396
rect 124236 4226 124516 4228
rect 124236 4174 124238 4226
rect 124290 4174 124516 4226
rect 124236 4172 124516 4174
rect 124236 4162 124292 4172
rect 123564 3614 123566 3666
rect 123618 3614 123620 3666
rect 123564 3602 123620 3614
rect 121436 3378 121492 3388
rect 121996 3444 122052 3454
rect 121996 3350 122052 3388
rect 122668 3444 122724 3454
rect 122780 3444 122836 3454
rect 122668 3442 122780 3444
rect 122668 3390 122670 3442
rect 122722 3390 122780 3442
rect 122668 3388 122780 3390
rect 122668 3378 122724 3388
rect 121324 1250 121380 1260
rect 122780 800 122836 3388
rect 124348 3444 124404 3454
rect 124348 3350 124404 3388
rect 124460 800 124516 4172
rect 124908 2996 124964 4956
rect 125132 5012 125188 5022
rect 125132 4918 125188 4956
rect 125916 4226 125972 5070
rect 126588 4340 126644 5740
rect 126812 5012 126868 5022
rect 126812 4918 126868 4956
rect 126924 4450 126980 8428
rect 127820 5794 127876 5806
rect 127820 5742 127822 5794
rect 127874 5742 127876 5794
rect 127596 5010 127652 5022
rect 127596 4958 127598 5010
rect 127650 4958 127652 5010
rect 127596 4676 127652 4958
rect 127596 4610 127652 4620
rect 126924 4398 126926 4450
rect 126978 4398 126980 4450
rect 126812 4340 126868 4350
rect 126588 4284 126812 4340
rect 125916 4174 125918 4226
rect 125970 4174 125972 4226
rect 126812 4208 126868 4284
rect 125916 4162 125972 4174
rect 126924 4116 126980 4398
rect 127820 4452 127876 5742
rect 127932 5010 127988 29260
rect 130082 29036 130346 29046
rect 130138 28980 130186 29036
rect 130242 28980 130290 29036
rect 130082 28970 130346 28980
rect 130082 27468 130346 27478
rect 130138 27412 130186 27468
rect 130242 27412 130290 27468
rect 130082 27402 130346 27412
rect 130082 25900 130346 25910
rect 130138 25844 130186 25900
rect 130242 25844 130290 25900
rect 130082 25834 130346 25844
rect 130082 24332 130346 24342
rect 130138 24276 130186 24332
rect 130242 24276 130290 24332
rect 130082 24266 130346 24276
rect 130082 22764 130346 22774
rect 130138 22708 130186 22764
rect 130242 22708 130290 22764
rect 130082 22698 130346 22708
rect 130082 21196 130346 21206
rect 130138 21140 130186 21196
rect 130242 21140 130290 21196
rect 130082 21130 130346 21140
rect 130082 19628 130346 19638
rect 130138 19572 130186 19628
rect 130242 19572 130290 19628
rect 130082 19562 130346 19572
rect 130082 18060 130346 18070
rect 130138 18004 130186 18060
rect 130242 18004 130290 18060
rect 130082 17994 130346 18004
rect 130082 16492 130346 16502
rect 130138 16436 130186 16492
rect 130242 16436 130290 16492
rect 130082 16426 130346 16436
rect 130082 14924 130346 14934
rect 130138 14868 130186 14924
rect 130242 14868 130290 14924
rect 130082 14858 130346 14868
rect 130508 14196 130564 14206
rect 130082 13356 130346 13366
rect 130138 13300 130186 13356
rect 130242 13300 130290 13356
rect 130082 13290 130346 13300
rect 130082 11788 130346 11798
rect 130138 11732 130186 11788
rect 130242 11732 130290 11788
rect 130082 11722 130346 11732
rect 130082 10220 130346 10230
rect 130138 10164 130186 10220
rect 130242 10164 130290 10220
rect 130082 10154 130346 10164
rect 130082 8652 130346 8662
rect 130138 8596 130186 8652
rect 130242 8596 130290 8652
rect 130082 8586 130346 8596
rect 129836 7588 129892 7598
rect 128828 6916 128884 6926
rect 128828 6690 128884 6860
rect 128828 6638 128830 6690
rect 128882 6638 128884 6690
rect 128828 6020 128884 6638
rect 129612 6692 129668 6702
rect 129836 6692 129892 7532
rect 130396 7362 130452 7374
rect 130396 7310 130398 7362
rect 130450 7310 130452 7362
rect 130396 7250 130452 7310
rect 130396 7198 130398 7250
rect 130450 7198 130452 7250
rect 130396 7186 130452 7198
rect 130082 7084 130346 7094
rect 130138 7028 130186 7084
rect 130242 7028 130290 7084
rect 130082 7018 130346 7028
rect 129612 6690 129892 6692
rect 129612 6638 129614 6690
rect 129666 6638 129892 6690
rect 129612 6636 129892 6638
rect 129612 6626 129668 6636
rect 130172 6580 130228 6590
rect 129724 6578 130228 6580
rect 129724 6526 130174 6578
rect 130226 6526 130228 6578
rect 129724 6524 130228 6526
rect 128828 5954 128884 5964
rect 129276 6466 129332 6478
rect 129276 6414 129278 6466
rect 129330 6414 129332 6466
rect 127932 4958 127934 5010
rect 127986 4958 127988 5010
rect 127932 4946 127988 4958
rect 128268 5794 128324 5806
rect 128268 5742 128270 5794
rect 128322 5742 128324 5794
rect 128268 5012 128324 5742
rect 128940 5796 128996 5806
rect 128940 5122 128996 5740
rect 128940 5070 128942 5122
rect 128994 5070 128996 5122
rect 128940 5058 128996 5070
rect 128828 5012 128884 5022
rect 128268 5010 128884 5012
rect 128268 4958 128830 5010
rect 128882 4958 128884 5010
rect 128268 4956 128884 4958
rect 127932 4676 127988 4686
rect 127932 4562 127988 4620
rect 127932 4510 127934 4562
rect 127986 4510 127988 4562
rect 127932 4498 127988 4510
rect 126476 4060 126980 4116
rect 127596 4116 127652 4126
rect 126476 3666 126532 4060
rect 127596 4022 127652 4060
rect 126476 3614 126478 3666
rect 126530 3614 126532 3666
rect 126476 3602 126532 3614
rect 126028 3444 126084 3454
rect 126140 3444 126196 3454
rect 126028 3442 126140 3444
rect 126028 3390 126030 3442
rect 126082 3390 126140 3442
rect 126028 3388 126140 3390
rect 126028 3378 126084 3388
rect 124908 2930 124964 2940
rect 126140 800 126196 3388
rect 127372 3444 127428 3454
rect 127372 3350 127428 3388
rect 127820 800 127876 4396
rect 128492 4116 128548 4126
rect 128492 3666 128548 4060
rect 128492 3614 128494 3666
rect 128546 3614 128548 3666
rect 128492 3602 128548 3614
rect 128828 1204 128884 4956
rect 129276 4564 129332 6414
rect 129500 6020 129556 6030
rect 129500 5926 129556 5964
rect 129724 5346 129780 6524
rect 130172 6514 130228 6524
rect 130508 6578 130564 14140
rect 130956 7588 131012 7598
rect 130844 7586 131012 7588
rect 130844 7534 130958 7586
rect 131010 7534 131012 7586
rect 130844 7532 131012 7534
rect 130508 6526 130510 6578
rect 130562 6526 130564 6578
rect 130508 6514 130564 6526
rect 130620 7250 130676 7262
rect 130620 7198 130622 7250
rect 130674 7198 130676 7250
rect 130508 6132 130564 6142
rect 130508 6038 130564 6076
rect 129948 6018 130004 6030
rect 129948 5966 129950 6018
rect 130002 5966 130004 6018
rect 129948 5796 130004 5966
rect 129948 5730 130004 5740
rect 130172 5684 130228 5694
rect 130172 5682 130564 5684
rect 130172 5630 130174 5682
rect 130226 5630 130564 5682
rect 130172 5628 130564 5630
rect 130172 5618 130228 5628
rect 130082 5516 130346 5526
rect 130138 5460 130186 5516
rect 130242 5460 130290 5516
rect 130082 5450 130346 5460
rect 129724 5294 129726 5346
rect 129778 5294 129780 5346
rect 129724 5282 129780 5294
rect 129276 4498 129332 4508
rect 129388 5122 129444 5134
rect 129388 5070 129390 5122
rect 129442 5070 129444 5122
rect 129164 4452 129220 4462
rect 129164 4358 129220 4396
rect 129276 4340 129332 4350
rect 129276 3668 129332 4284
rect 129388 4228 129444 5070
rect 130284 4228 130340 4238
rect 129388 4226 130340 4228
rect 129388 4174 130286 4226
rect 130338 4174 130340 4226
rect 129388 4172 130340 4174
rect 130284 4162 130340 4172
rect 130082 3948 130346 3958
rect 130138 3892 130186 3948
rect 130242 3892 130290 3948
rect 130082 3882 130346 3892
rect 129276 3536 129332 3612
rect 129836 3668 129892 3678
rect 129836 3574 129892 3612
rect 130508 3668 130564 5628
rect 130620 5010 130676 7198
rect 130620 4958 130622 5010
rect 130674 4958 130676 5010
rect 130620 4788 130676 4958
rect 130620 4722 130676 4732
rect 130844 5012 130900 7532
rect 130956 7522 131012 7532
rect 131292 7588 131348 7598
rect 131292 7494 131348 7532
rect 131068 6578 131124 6590
rect 131068 6526 131070 6578
rect 131122 6526 131124 6578
rect 131068 6132 131124 6526
rect 131404 6578 131460 30828
rect 131964 11956 132020 11966
rect 131740 7588 131796 7598
rect 131740 7494 131796 7532
rect 131404 6526 131406 6578
rect 131458 6526 131460 6578
rect 131404 6514 131460 6526
rect 131964 6690 132020 11900
rect 131964 6638 131966 6690
rect 132018 6638 132020 6690
rect 131068 6066 131124 6076
rect 131740 6020 131796 6030
rect 131964 6020 132020 6638
rect 132972 6578 133028 6590
rect 132972 6526 132974 6578
rect 133026 6526 133028 6578
rect 131740 6018 132020 6020
rect 131740 5966 131742 6018
rect 131794 5966 132020 6018
rect 131740 5964 132020 5966
rect 132076 6018 132132 6030
rect 132076 5966 132078 6018
rect 132130 5966 132132 6018
rect 131740 5954 131796 5964
rect 130956 5796 131012 5806
rect 130956 5122 131012 5740
rect 132076 5796 132132 5966
rect 132636 5908 132692 5918
rect 132636 5814 132692 5852
rect 132076 5730 132132 5740
rect 132300 5682 132356 5694
rect 132300 5630 132302 5682
rect 132354 5630 132356 5682
rect 131740 5348 131796 5358
rect 131740 5254 131796 5292
rect 130956 5070 130958 5122
rect 131010 5070 131012 5122
rect 130956 5058 131012 5070
rect 131404 5122 131460 5134
rect 131404 5070 131406 5122
rect 131458 5070 131460 5122
rect 130508 3602 130564 3612
rect 129500 3556 129556 3566
rect 128828 1138 128884 1148
rect 129500 800 129556 3500
rect 130396 3444 130452 3454
rect 130844 3444 130900 4956
rect 131404 4226 131460 5070
rect 131404 4174 131406 4226
rect 131458 4174 131460 4226
rect 131404 4162 131460 4174
rect 132300 4228 132356 5630
rect 132972 5348 133028 6526
rect 133308 6578 133364 31500
rect 133532 12068 133588 12078
rect 133532 7700 133588 12012
rect 133532 7634 133588 7644
rect 133980 10388 134036 10398
rect 133308 6526 133310 6578
rect 133362 6526 133364 6578
rect 133308 6514 133364 6526
rect 133644 6468 133700 6478
rect 132972 5282 133028 5292
rect 133308 5906 133364 5918
rect 133308 5854 133310 5906
rect 133362 5854 133364 5906
rect 132972 5012 133028 5022
rect 132972 4918 133028 4956
rect 133308 5012 133364 5854
rect 133532 5124 133588 5134
rect 133532 5030 133588 5068
rect 132300 4162 132356 4172
rect 132412 4450 132468 4462
rect 132412 4398 132414 4450
rect 132466 4398 132468 4450
rect 131180 3668 131236 3678
rect 131180 3574 131236 3612
rect 132188 3556 132244 3566
rect 130396 3442 130900 3444
rect 130396 3390 130398 3442
rect 130450 3390 130900 3442
rect 130396 3388 130900 3390
rect 131180 3444 131236 3454
rect 130396 3378 130452 3388
rect 131180 800 131236 3388
rect 132188 3442 132244 3500
rect 132188 3390 132190 3442
rect 132242 3390 132244 3442
rect 132188 3378 132244 3390
rect 132412 3444 132468 4398
rect 132412 3378 132468 3388
rect 132860 4452 132916 4462
rect 132860 800 132916 4396
rect 133308 3554 133364 4956
rect 133420 4228 133476 4238
rect 133420 4134 133476 4172
rect 133644 3892 133700 6412
rect 133980 6466 134036 10332
rect 133980 6414 133982 6466
rect 134034 6414 134036 6466
rect 133756 5796 133812 5806
rect 133756 5702 133812 5740
rect 133980 5684 134036 6414
rect 134764 6130 134820 33068
rect 134764 6078 134766 6130
rect 134818 6078 134820 6130
rect 134764 6066 134820 6078
rect 136220 8820 136276 8830
rect 136220 6132 136276 8764
rect 137004 6468 137060 6478
rect 137004 6374 137060 6412
rect 136220 6000 136276 6076
rect 137340 6130 137396 33964
rect 138572 29988 138628 29998
rect 138572 14196 138628 29932
rect 138572 14130 138628 14140
rect 137564 10500 137620 10510
rect 137564 6690 137620 10444
rect 139020 7698 139076 36204
rect 142156 36260 142212 36270
rect 142156 36166 142212 36204
rect 143052 36260 143108 36430
rect 144844 36482 144900 36494
rect 144844 36430 144846 36482
rect 144898 36430 144900 36482
rect 143052 36194 143108 36204
rect 144172 36372 144228 36382
rect 142156 35588 142212 35598
rect 141260 34692 141316 34702
rect 141036 28644 141092 28654
rect 139468 23044 139524 23054
rect 139468 14420 139524 22988
rect 141036 22932 141092 28588
rect 141036 22866 141092 22876
rect 139468 14354 139524 14364
rect 140028 12404 140084 12414
rect 139020 7646 139022 7698
rect 139074 7646 139076 7698
rect 139020 7634 139076 7646
rect 139916 7700 139972 7710
rect 139916 7606 139972 7644
rect 138796 7476 138852 7486
rect 138796 7474 139300 7476
rect 138796 7422 138798 7474
rect 138850 7422 139300 7474
rect 138796 7420 139300 7422
rect 138796 7410 138852 7420
rect 137564 6638 137566 6690
rect 137618 6638 137620 6690
rect 137564 6580 137620 6638
rect 137564 6514 137620 6524
rect 137788 7362 137844 7374
rect 137788 7310 137790 7362
rect 137842 7310 137844 7362
rect 137788 6468 137844 7310
rect 139244 6914 139300 7420
rect 139244 6862 139246 6914
rect 139298 6862 139300 6914
rect 139244 6850 139300 6862
rect 139692 7474 139748 7486
rect 139692 7422 139694 7474
rect 139746 7422 139748 7474
rect 138908 6802 138964 6814
rect 138908 6750 138910 6802
rect 138962 6750 138964 6802
rect 138124 6580 138180 6590
rect 138124 6486 138180 6524
rect 138684 6578 138740 6590
rect 138684 6526 138686 6578
rect 138738 6526 138740 6578
rect 137788 6402 137844 6412
rect 138684 6468 138740 6526
rect 138908 6580 138964 6750
rect 138908 6514 138964 6524
rect 137340 6078 137342 6130
rect 137394 6078 137396 6130
rect 137340 6066 137396 6078
rect 138236 6132 138292 6142
rect 138236 6018 138292 6076
rect 138236 5966 138238 6018
rect 138290 5966 138292 6018
rect 138236 5954 138292 5966
rect 138684 6020 138740 6412
rect 139692 6132 139748 7422
rect 139916 6692 139972 6702
rect 140028 6692 140084 12348
rect 140364 7362 140420 7374
rect 140364 7310 140366 7362
rect 140418 7310 140420 7362
rect 139916 6690 140196 6692
rect 139916 6638 139918 6690
rect 139970 6638 140196 6690
rect 139916 6636 140196 6638
rect 139916 6626 139972 6636
rect 139692 6066 139748 6076
rect 138684 5926 138740 5964
rect 140140 6018 140196 6636
rect 140140 5966 140142 6018
rect 140194 5966 140196 6018
rect 140140 5954 140196 5966
rect 140364 6020 140420 7310
rect 134428 5908 134484 5918
rect 134428 5814 134484 5852
rect 137004 5906 137060 5918
rect 137004 5854 137006 5906
rect 137058 5854 137060 5906
rect 135884 5794 135940 5806
rect 135884 5742 135886 5794
rect 135938 5742 135940 5794
rect 133980 5628 134484 5684
rect 134428 5010 134484 5628
rect 135436 5348 135492 5358
rect 135436 5254 135492 5292
rect 134652 5124 134708 5134
rect 134652 5030 134708 5068
rect 135100 5122 135156 5134
rect 135100 5070 135102 5122
rect 135154 5070 135156 5122
rect 134428 4958 134430 5010
rect 134482 4958 134484 5010
rect 134428 4946 134484 4958
rect 134428 4452 134484 4462
rect 134428 4358 134484 4396
rect 133644 3666 133700 3836
rect 133644 3614 133646 3666
rect 133698 3614 133700 3666
rect 133644 3602 133700 3614
rect 135100 3666 135156 5070
rect 135884 5012 135940 5742
rect 137004 5348 137060 5854
rect 140364 5906 140420 5964
rect 140364 5854 140366 5906
rect 140418 5854 140420 5906
rect 140364 5842 140420 5854
rect 140924 6578 140980 6590
rect 140924 6526 140926 6578
rect 140978 6526 140980 6578
rect 138908 5684 138964 5694
rect 139244 5684 139300 5694
rect 138908 5590 138964 5628
rect 139020 5682 139300 5684
rect 139020 5630 139246 5682
rect 139298 5630 139300 5682
rect 139020 5628 139300 5630
rect 137004 5282 137060 5292
rect 137340 5460 137396 5470
rect 137340 5346 137396 5404
rect 139020 5348 139076 5628
rect 139244 5618 139300 5628
rect 140812 5682 140868 5694
rect 140812 5630 140814 5682
rect 140866 5630 140868 5682
rect 137340 5294 137342 5346
rect 137394 5294 137396 5346
rect 137340 5282 137396 5294
rect 137900 5292 139076 5348
rect 139244 5348 139300 5358
rect 136556 5124 136612 5134
rect 136556 5030 136612 5068
rect 137004 5122 137060 5134
rect 137004 5070 137006 5122
rect 137058 5070 137060 5122
rect 135884 4946 135940 4956
rect 136444 5012 136500 5022
rect 135772 4452 135828 4462
rect 135772 4358 135828 4396
rect 135100 3614 135102 3666
rect 135154 3614 135156 3666
rect 135100 3602 135156 3614
rect 135324 4226 135380 4238
rect 136220 4228 136276 4238
rect 135324 4174 135326 4226
rect 135378 4174 135380 4226
rect 133308 3502 133310 3554
rect 133362 3502 133364 3554
rect 133308 3490 133364 3502
rect 135324 3556 135380 4174
rect 135324 3490 135380 3500
rect 136108 4226 136276 4228
rect 136108 4174 136222 4226
rect 136274 4174 136276 4226
rect 136108 4172 136276 4174
rect 134204 3444 134260 3454
rect 134204 3350 134260 3388
rect 134540 3444 134596 3454
rect 134540 800 134596 3388
rect 136108 3444 136164 4172
rect 136220 4162 136276 4172
rect 136108 3350 136164 3388
rect 136220 3556 136276 3566
rect 136220 800 136276 3500
rect 136444 980 136500 4956
rect 137004 4226 137060 5070
rect 137004 4174 137006 4226
rect 137058 4174 137060 4226
rect 137004 4162 137060 4174
rect 137004 3556 137060 3566
rect 137004 3462 137060 3500
rect 137900 3554 137956 5292
rect 139244 5254 139300 5292
rect 138460 5124 138516 5134
rect 138460 5030 138516 5068
rect 138908 5122 138964 5134
rect 138908 5070 138910 5122
rect 138962 5070 138964 5122
rect 138348 5012 138404 5022
rect 137900 3502 137902 3554
rect 137954 3502 137956 3554
rect 137900 3490 137956 3502
rect 138012 4450 138068 4462
rect 138012 4398 138014 4450
rect 138066 4398 138068 4450
rect 138012 3444 138068 4398
rect 138012 3378 138068 3388
rect 138124 4228 138180 4238
rect 138124 2884 138180 4172
rect 138236 3332 138292 3342
rect 138236 3238 138292 3276
rect 136444 914 136500 924
rect 137900 2828 138180 2884
rect 137900 800 137956 2828
rect 138348 1428 138404 4956
rect 138908 3668 138964 5070
rect 139804 5122 139860 5134
rect 139804 5070 139806 5122
rect 139858 5070 139860 5122
rect 139804 5012 139860 5070
rect 139804 4946 139860 4956
rect 140140 4450 140196 4462
rect 140140 4398 140142 4450
rect 140194 4398 140196 4450
rect 139020 4228 139076 4238
rect 139020 4134 139076 4172
rect 140028 4228 140084 4238
rect 139020 3668 139076 3678
rect 138908 3666 139076 3668
rect 138908 3614 139022 3666
rect 139074 3614 139076 3666
rect 138908 3612 139076 3614
rect 139020 3602 139076 3612
rect 138348 1362 138404 1372
rect 139580 3444 139636 3454
rect 139580 800 139636 3388
rect 140028 3442 140084 4172
rect 140028 3390 140030 3442
rect 140082 3390 140084 3442
rect 140028 3378 140084 3390
rect 140140 3444 140196 4398
rect 140812 4228 140868 5630
rect 140924 5460 140980 6526
rect 141260 6578 141316 34636
rect 141260 6526 141262 6578
rect 141314 6526 141316 6578
rect 141260 6514 141316 6526
rect 141148 6132 141204 6142
rect 141148 6038 141204 6076
rect 142156 6130 142212 35532
rect 143836 35588 143892 35598
rect 144172 35588 144228 36316
rect 144844 36372 144900 36430
rect 147084 36482 147140 36494
rect 147084 36430 147086 36482
rect 147138 36430 147140 36482
rect 144844 36306 144900 36316
rect 145964 36370 146020 36382
rect 145964 36318 145966 36370
rect 146018 36318 146020 36370
rect 145964 36260 146020 36318
rect 145964 36194 146020 36204
rect 144956 35698 145012 35710
rect 146748 35700 146804 35710
rect 144956 35646 144958 35698
rect 145010 35646 145012 35698
rect 143836 35586 144228 35588
rect 143836 35534 143838 35586
rect 143890 35534 144228 35586
rect 143836 35532 144228 35534
rect 143836 35522 143892 35532
rect 143500 21476 143556 21486
rect 142716 9604 142772 9614
rect 142716 8428 142772 9548
rect 142716 8372 142996 8428
rect 142156 6078 142158 6130
rect 142210 6078 142212 6130
rect 142156 6066 142212 6078
rect 142716 8036 142772 8046
rect 140924 5394 140980 5404
rect 141820 5906 141876 5918
rect 141820 5854 141822 5906
rect 141874 5854 141876 5906
rect 141820 5348 141876 5854
rect 142716 5794 142772 7980
rect 142940 6802 142996 8372
rect 142940 6750 142942 6802
rect 142994 6750 142996 6802
rect 142940 6738 142996 6750
rect 142716 5742 142718 5794
rect 142770 5742 142772 5794
rect 142716 5730 142772 5742
rect 143164 6580 143220 6590
rect 141820 5282 141876 5292
rect 142940 5684 142996 5694
rect 142940 5234 142996 5628
rect 142940 5182 142942 5234
rect 142994 5182 142996 5234
rect 142940 5170 142996 5182
rect 141148 5124 141204 5134
rect 141820 5124 141876 5134
rect 141148 5030 141204 5068
rect 141596 5122 141876 5124
rect 141596 5070 141822 5122
rect 141874 5070 141876 5122
rect 141596 5068 141876 5070
rect 141260 5010 141316 5022
rect 141260 4958 141262 5010
rect 141314 4958 141316 5010
rect 141260 4900 141316 4958
rect 140812 4162 140868 4172
rect 141148 4844 141316 4900
rect 141148 3780 141204 4844
rect 141260 4228 141316 4238
rect 141596 4228 141652 5068
rect 141820 5058 141876 5068
rect 142156 4898 142212 4910
rect 142156 4846 142158 4898
rect 142210 4846 142212 4898
rect 142156 4452 142212 4846
rect 142828 4452 142884 4462
rect 142156 4386 142212 4396
rect 142716 4450 142884 4452
rect 142716 4398 142830 4450
rect 142882 4398 142884 4450
rect 142716 4396 142884 4398
rect 141260 4226 141652 4228
rect 141260 4174 141262 4226
rect 141314 4174 141652 4226
rect 141260 4172 141652 4174
rect 141820 4228 141876 4238
rect 141260 4162 141316 4172
rect 141820 4134 141876 4172
rect 142044 4228 142100 4238
rect 141148 3714 141204 3724
rect 141484 3780 141540 3790
rect 141484 3666 141540 3724
rect 141484 3614 141486 3666
rect 141538 3614 141540 3666
rect 141484 3602 141540 3614
rect 140140 3378 140196 3388
rect 140924 3444 140980 3454
rect 140924 3350 140980 3388
rect 141260 3444 141316 3454
rect 141260 800 141316 3388
rect 141820 3444 141876 3454
rect 141820 3350 141876 3388
rect 142044 2660 142100 4172
rect 142716 3444 142772 4396
rect 142828 4386 142884 4396
rect 143164 3666 143220 6524
rect 143500 5908 143556 21420
rect 143500 5842 143556 5852
rect 143948 19012 144004 19022
rect 143836 4452 143892 4462
rect 143836 4358 143892 4396
rect 143164 3614 143166 3666
rect 143218 3614 143220 3666
rect 143164 3602 143220 3614
rect 142716 3378 142772 3388
rect 142940 3444 142996 3454
rect 142044 2594 142100 2604
rect 142940 800 142996 3388
rect 143948 2548 144004 18956
rect 144060 6018 144116 6030
rect 144060 5966 144062 6018
rect 144114 5966 144116 6018
rect 144060 5796 144116 5966
rect 144060 5730 144116 5740
rect 144172 4562 144228 35532
rect 144284 35588 144340 35598
rect 144284 35494 144340 35532
rect 144956 35588 145012 35646
rect 146636 35698 146804 35700
rect 146636 35646 146750 35698
rect 146802 35646 146804 35698
rect 146636 35644 146804 35646
rect 144956 35522 145012 35532
rect 146076 35586 146132 35598
rect 146076 35534 146078 35586
rect 146130 35534 146132 35586
rect 146076 35252 146132 35534
rect 146076 35186 146132 35196
rect 144956 34914 145012 34926
rect 144956 34862 144958 34914
rect 145010 34862 145012 34914
rect 144396 34692 144452 34702
rect 144396 34598 144452 34636
rect 144956 34692 145012 34862
rect 144956 34626 145012 34636
rect 146076 34802 146132 34814
rect 146076 34750 146078 34802
rect 146130 34750 146132 34802
rect 146076 34356 146132 34750
rect 146636 34692 146692 35644
rect 146748 35634 146804 35644
rect 146636 34598 146692 34636
rect 147084 34690 147140 36430
rect 147644 35586 147700 38780
rect 147756 37044 147812 37054
rect 147756 36594 147812 36988
rect 147756 36542 147758 36594
rect 147810 36542 147812 36594
rect 147756 36530 147812 36542
rect 148492 36092 148756 36102
rect 148548 36036 148596 36092
rect 148652 36036 148700 36092
rect 148492 36026 148756 36036
rect 147644 35534 147646 35586
rect 147698 35534 147700 35586
rect 147644 35522 147700 35534
rect 147084 34638 147086 34690
rect 147138 34638 147140 34690
rect 146076 34290 146132 34300
rect 144956 34130 145012 34142
rect 144956 34078 144958 34130
rect 145010 34078 145012 34130
rect 144284 34020 144340 34030
rect 144284 33926 144340 33964
rect 144956 34020 145012 34078
rect 144956 33954 145012 33964
rect 146076 34018 146132 34030
rect 146076 33966 146078 34018
rect 146130 33966 146132 34018
rect 146076 33460 146132 33966
rect 146076 33394 146132 33404
rect 144956 33346 145012 33358
rect 144956 33294 144958 33346
rect 145010 33294 145012 33346
rect 144396 33124 144452 33134
rect 144396 33030 144452 33068
rect 144956 33124 145012 33294
rect 144956 33058 145012 33068
rect 146076 33234 146132 33246
rect 146076 33182 146078 33234
rect 146130 33182 146132 33234
rect 146076 32564 146132 33182
rect 146076 32498 146132 32508
rect 144956 31778 145012 31790
rect 144956 31726 144958 31778
rect 145010 31726 145012 31778
rect 144396 31556 144452 31566
rect 144396 31462 144452 31500
rect 144956 31556 145012 31726
rect 146076 31668 146132 31678
rect 146076 31574 146132 31612
rect 144956 31490 145012 31500
rect 144956 30994 145012 31006
rect 144956 30942 144958 30994
rect 145010 30942 145012 30994
rect 144284 30884 144340 30894
rect 144284 30790 144340 30828
rect 144956 30884 145012 30942
rect 144956 30818 145012 30828
rect 146076 30882 146132 30894
rect 146076 30830 146078 30882
rect 146130 30830 146132 30882
rect 146076 30772 146132 30830
rect 146076 30706 146132 30716
rect 144956 30210 145012 30222
rect 144956 30158 144958 30210
rect 145010 30158 145012 30210
rect 144396 29988 144452 29998
rect 144396 29894 144452 29932
rect 144956 29988 145012 30158
rect 144956 29922 145012 29932
rect 146076 30098 146132 30110
rect 146076 30046 146078 30098
rect 146130 30046 146132 30098
rect 146076 29988 146132 30046
rect 146076 29922 146132 29932
rect 144956 29426 145012 29438
rect 144956 29374 144958 29426
rect 145010 29374 145012 29426
rect 144284 29316 144340 29326
rect 144284 29222 144340 29260
rect 144956 29316 145012 29374
rect 144956 29250 145012 29260
rect 146076 29314 146132 29326
rect 146076 29262 146078 29314
rect 146130 29262 146132 29314
rect 146076 28980 146132 29262
rect 146076 28914 146132 28924
rect 144396 28644 144452 28654
rect 144396 28550 144452 28588
rect 144956 28644 145012 28654
rect 144956 28550 145012 28588
rect 146076 28642 146132 28654
rect 146076 28590 146078 28642
rect 146130 28590 146132 28642
rect 146076 28084 146132 28590
rect 146076 28018 146132 28028
rect 144956 27858 145012 27870
rect 144956 27806 144958 27858
rect 145010 27806 145012 27858
rect 144284 27748 144340 27758
rect 144284 27654 144340 27692
rect 144956 27748 145012 27806
rect 144956 27682 145012 27692
rect 146076 27746 146132 27758
rect 146076 27694 146078 27746
rect 146130 27694 146132 27746
rect 146076 27188 146132 27694
rect 146076 27122 146132 27132
rect 144956 27074 145012 27086
rect 144956 27022 144958 27074
rect 145010 27022 145012 27074
rect 144396 26964 144452 26974
rect 144396 26870 144452 26908
rect 144956 26964 145012 27022
rect 144956 26898 145012 26908
rect 146076 26962 146132 26974
rect 146076 26910 146078 26962
rect 146130 26910 146132 26962
rect 146076 26292 146132 26910
rect 146076 26226 146132 26236
rect 144956 25506 145012 25518
rect 144956 25454 144958 25506
rect 145010 25454 145012 25506
rect 144396 25284 144452 25294
rect 144396 25190 144452 25228
rect 144956 25284 145012 25454
rect 146076 25396 146132 25406
rect 146076 25302 146132 25340
rect 144956 25218 145012 25228
rect 144956 24722 145012 24734
rect 144956 24670 144958 24722
rect 145010 24670 145012 24722
rect 144284 24612 144340 24622
rect 144284 24518 144340 24556
rect 144956 24612 145012 24670
rect 144956 24546 145012 24556
rect 146076 24610 146132 24622
rect 146076 24558 146078 24610
rect 146130 24558 146132 24610
rect 146076 24500 146132 24558
rect 146076 24434 146132 24444
rect 144956 23938 145012 23950
rect 144956 23886 144958 23938
rect 145010 23886 145012 23938
rect 144396 23716 144452 23726
rect 144396 23622 144452 23660
rect 144956 23716 145012 23886
rect 144956 23650 145012 23660
rect 146076 23826 146132 23838
rect 146076 23774 146078 23826
rect 146130 23774 146132 23826
rect 146076 23716 146132 23774
rect 146076 23650 146132 23660
rect 144956 23154 145012 23166
rect 144956 23102 144958 23154
rect 145010 23102 145012 23154
rect 144284 23044 144340 23054
rect 144284 22950 144340 22988
rect 144956 23044 145012 23102
rect 144956 22978 145012 22988
rect 146076 23042 146132 23054
rect 146076 22990 146078 23042
rect 146130 22990 146132 23042
rect 146076 22708 146132 22990
rect 146076 22642 146132 22652
rect 144956 22370 145012 22382
rect 144956 22318 144958 22370
rect 145010 22318 145012 22370
rect 144396 22148 144452 22158
rect 144396 22054 144452 22092
rect 144956 22148 145012 22318
rect 144956 22082 145012 22092
rect 146076 22258 146132 22270
rect 146076 22206 146078 22258
rect 146130 22206 146132 22258
rect 146076 21812 146132 22206
rect 146076 21746 146132 21756
rect 144956 21586 145012 21598
rect 144956 21534 144958 21586
rect 145010 21534 145012 21586
rect 144284 21476 144340 21486
rect 144284 21382 144340 21420
rect 144956 21476 145012 21534
rect 144956 21410 145012 21420
rect 146076 21474 146132 21486
rect 146076 21422 146078 21474
rect 146130 21422 146132 21474
rect 146076 20916 146132 21422
rect 146076 20850 146132 20860
rect 144956 20802 145012 20814
rect 144956 20750 144958 20802
rect 145010 20750 145012 20802
rect 144396 20580 144452 20590
rect 144396 20486 144452 20524
rect 144956 20580 145012 20750
rect 144956 20514 145012 20524
rect 146076 20690 146132 20702
rect 146076 20638 146078 20690
rect 146130 20638 146132 20690
rect 146076 20020 146132 20638
rect 146076 19954 146132 19964
rect 144956 19234 145012 19246
rect 144956 19182 144958 19234
rect 145010 19182 145012 19234
rect 144396 19012 144452 19022
rect 144396 18918 144452 18956
rect 144956 19012 145012 19182
rect 146076 19124 146132 19134
rect 146076 19030 146132 19068
rect 144956 18946 145012 18956
rect 144956 18450 145012 18462
rect 144956 18398 144958 18450
rect 145010 18398 145012 18450
rect 144284 18340 144340 18350
rect 144284 18246 144340 18284
rect 144956 18340 145012 18398
rect 144956 18274 145012 18284
rect 146076 18338 146132 18350
rect 146076 18286 146078 18338
rect 146130 18286 146132 18338
rect 146076 18228 146132 18286
rect 146076 18162 146132 18172
rect 144956 17666 145012 17678
rect 144956 17614 144958 17666
rect 145010 17614 145012 17666
rect 144396 17444 144452 17454
rect 144396 17350 144452 17388
rect 144956 17444 145012 17614
rect 144956 17378 145012 17388
rect 146076 17554 146132 17566
rect 146076 17502 146078 17554
rect 146130 17502 146132 17554
rect 146076 17444 146132 17502
rect 146076 17378 146132 17388
rect 144284 16884 144340 16894
rect 144284 16790 144340 16828
rect 144956 16884 145012 16894
rect 144956 16790 145012 16828
rect 146076 16882 146132 16894
rect 146076 16830 146078 16882
rect 146130 16830 146132 16882
rect 146076 16436 146132 16830
rect 146076 16370 146132 16380
rect 144956 16098 145012 16110
rect 144956 16046 144958 16098
rect 145010 16046 145012 16098
rect 144396 15876 144452 15886
rect 144396 15782 144452 15820
rect 144956 15876 145012 16046
rect 144956 15810 145012 15820
rect 146076 15986 146132 15998
rect 146076 15934 146078 15986
rect 146130 15934 146132 15986
rect 146076 15540 146132 15934
rect 146076 15474 146132 15484
rect 144284 15316 144340 15326
rect 144284 15202 144340 15260
rect 144956 15316 145012 15326
rect 144956 15222 145012 15260
rect 144284 15150 144286 15202
rect 144338 15150 144340 15202
rect 144284 12852 144340 15150
rect 146076 15202 146132 15214
rect 146076 15150 146078 15202
rect 146130 15150 146132 15202
rect 146076 14644 146132 15150
rect 146076 14578 146132 14588
rect 144956 14530 145012 14542
rect 144956 14478 144958 14530
rect 145010 14478 145012 14530
rect 144396 14308 144452 14318
rect 144396 14214 144452 14252
rect 144956 14308 145012 14478
rect 144956 14242 145012 14252
rect 146076 14418 146132 14430
rect 146076 14366 146078 14418
rect 146130 14366 146132 14418
rect 146076 13748 146132 14366
rect 146076 13682 146132 13692
rect 144284 12786 144340 12796
rect 144396 12964 144452 12974
rect 144396 12738 144452 12908
rect 144956 12964 145012 12974
rect 144956 12870 145012 12908
rect 146076 12852 146132 12862
rect 146076 12758 146132 12796
rect 144396 12686 144398 12738
rect 144450 12686 144452 12738
rect 144284 12068 144340 12078
rect 144284 11974 144340 12012
rect 144396 11844 144452 12686
rect 144284 11788 144452 11844
rect 144620 12292 144676 12302
rect 144284 11172 144340 11788
rect 144284 11106 144340 11116
rect 144396 11170 144452 11182
rect 144396 11118 144398 11170
rect 144450 11118 144452 11170
rect 144396 10836 144452 11118
rect 144396 10770 144452 10780
rect 144284 7362 144340 7374
rect 144284 7310 144286 7362
rect 144338 7310 144340 7362
rect 144284 6580 144340 7310
rect 144284 6486 144340 6524
rect 144620 5236 144676 12236
rect 144956 12178 145012 12190
rect 144956 12126 144958 12178
rect 145010 12126 145012 12178
rect 144956 12068 145012 12126
rect 144956 12002 145012 12012
rect 146076 12066 146132 12078
rect 146076 12014 146078 12066
rect 146130 12014 146132 12066
rect 146076 11956 146132 12014
rect 146076 11890 146132 11900
rect 144956 11394 145012 11406
rect 144956 11342 144958 11394
rect 145010 11342 145012 11394
rect 144956 10836 145012 11342
rect 146076 11282 146132 11294
rect 146076 11230 146078 11282
rect 146130 11230 146132 11282
rect 146076 11172 146132 11230
rect 146076 11106 146132 11116
rect 144956 10770 145012 10780
rect 146300 10722 146356 10734
rect 146300 10670 146302 10722
rect 146354 10670 146356 10722
rect 145180 10498 145236 10510
rect 145180 10446 145182 10498
rect 145234 10446 145236 10498
rect 144956 9940 145012 9950
rect 144956 9846 145012 9884
rect 144956 8932 145012 8942
rect 144956 8838 145012 8876
rect 144956 8370 145012 8382
rect 144956 8318 144958 8370
rect 145010 8318 145012 8370
rect 144956 7924 145012 8318
rect 144732 7868 145012 7924
rect 144732 6692 144788 7868
rect 145068 7812 145124 7822
rect 144956 7476 145012 7486
rect 144956 7362 145012 7420
rect 144956 7310 144958 7362
rect 145010 7310 145012 7362
rect 144956 7298 145012 7310
rect 145068 6802 145124 7756
rect 145180 7588 145236 10446
rect 146300 10164 146356 10670
rect 146300 10098 146356 10108
rect 146860 10498 146916 10510
rect 146860 10446 146862 10498
rect 146914 10446 146916 10498
rect 146860 10164 146916 10446
rect 146860 10098 146916 10108
rect 146300 9716 146356 9726
rect 146300 9622 146356 9660
rect 146972 9716 147028 9726
rect 146972 9602 147028 9660
rect 146972 9550 146974 9602
rect 147026 9550 147028 9602
rect 146972 9268 147028 9550
rect 146972 9202 147028 9212
rect 146300 9156 146356 9166
rect 146300 9062 146356 9100
rect 146860 9156 146916 9166
rect 146860 8930 146916 9100
rect 146860 8878 146862 8930
rect 146914 8878 146916 8930
rect 146860 8484 146916 8878
rect 146860 8418 146916 8428
rect 146300 8148 146356 8158
rect 146300 8054 146356 8092
rect 146972 8148 147028 8158
rect 146972 8034 147028 8092
rect 146972 7982 146974 8034
rect 147026 7982 147028 8034
rect 146188 7588 146244 7598
rect 145180 7522 145236 7532
rect 146076 7532 146188 7588
rect 145068 6750 145070 6802
rect 145122 6750 145124 6802
rect 145068 6738 145124 6750
rect 144732 6626 144788 6636
rect 145180 6580 145236 6590
rect 144956 6244 145012 6254
rect 144956 5794 145012 6188
rect 144956 5742 144958 5794
rect 145010 5742 145012 5794
rect 144956 5730 145012 5742
rect 144956 5236 145012 5246
rect 144620 5234 145012 5236
rect 144620 5182 144958 5234
rect 145010 5182 145012 5234
rect 144620 5180 145012 5182
rect 144956 5170 145012 5180
rect 144284 5012 144340 5022
rect 144620 5012 144676 5022
rect 144284 5010 144620 5012
rect 144284 4958 144286 5010
rect 144338 4958 144620 5010
rect 144284 4956 144620 4958
rect 144284 4946 144340 4956
rect 144172 4510 144174 4562
rect 144226 4510 144228 4562
rect 144172 4498 144228 4510
rect 144172 3444 144228 3454
rect 144172 3350 144228 3388
rect 143948 2482 144004 2492
rect 144620 800 144676 4956
rect 144956 4228 145012 4238
rect 144956 4134 145012 4172
rect 145068 3444 145124 3454
rect 145068 3350 145124 3388
rect 145180 2996 145236 6524
rect 145180 2930 145236 2940
rect 145964 5796 146020 5806
rect 145964 1204 146020 5740
rect 146076 2100 146132 7532
rect 146188 7456 146244 7532
rect 146860 7588 146916 7598
rect 146860 7494 146916 7532
rect 146972 7476 147028 7982
rect 147084 7700 147140 34638
rect 147084 7634 147140 7644
rect 147868 34692 147924 34702
rect 146972 7410 147028 7420
rect 146300 6580 146356 6590
rect 146300 6486 146356 6524
rect 146972 6580 147028 6590
rect 146972 6486 147028 6524
rect 146300 6018 146356 6030
rect 146300 5966 146302 6018
rect 146354 5966 146356 6018
rect 146300 5684 146356 5966
rect 146860 5796 146916 5806
rect 146860 5702 146916 5740
rect 147308 5794 147364 5806
rect 147308 5742 147310 5794
rect 147362 5742 147364 5794
rect 146300 5618 146356 5628
rect 147308 5684 147364 5742
rect 147308 5618 147364 5628
rect 146860 5122 146916 5134
rect 146860 5070 146862 5122
rect 146914 5070 146916 5122
rect 146300 5010 146356 5022
rect 146300 4958 146302 5010
rect 146354 4958 146356 5010
rect 146300 4900 146356 4958
rect 146860 5012 146916 5070
rect 146860 4946 146916 4956
rect 146300 4834 146356 4844
rect 147420 4900 147476 4910
rect 147420 4806 147476 4844
rect 146300 4450 146356 4462
rect 146300 4398 146302 4450
rect 146354 4398 146356 4450
rect 146300 3892 146356 4398
rect 146300 3826 146356 3836
rect 146860 4226 146916 4238
rect 146860 4174 146862 4226
rect 146914 4174 146916 4226
rect 146860 3892 146916 4174
rect 146860 3826 146916 3836
rect 147868 3332 147924 34636
rect 148492 34524 148756 34534
rect 148548 34468 148596 34524
rect 148652 34468 148700 34524
rect 148492 34458 148756 34468
rect 148492 32956 148756 32966
rect 148548 32900 148596 32956
rect 148652 32900 148700 32956
rect 148492 32890 148756 32900
rect 148492 31388 148756 31398
rect 148548 31332 148596 31388
rect 148652 31332 148700 31388
rect 148492 31322 148756 31332
rect 148492 29820 148756 29830
rect 148548 29764 148596 29820
rect 148652 29764 148700 29820
rect 148492 29754 148756 29764
rect 148492 28252 148756 28262
rect 148548 28196 148596 28252
rect 148652 28196 148700 28252
rect 148492 28186 148756 28196
rect 148492 26684 148756 26694
rect 148548 26628 148596 26684
rect 148652 26628 148700 26684
rect 148492 26618 148756 26628
rect 148492 25116 148756 25126
rect 148548 25060 148596 25116
rect 148652 25060 148700 25116
rect 148492 25050 148756 25060
rect 148492 23548 148756 23558
rect 148548 23492 148596 23548
rect 148652 23492 148700 23548
rect 148492 23482 148756 23492
rect 148492 21980 148756 21990
rect 148548 21924 148596 21980
rect 148652 21924 148700 21980
rect 148492 21914 148756 21924
rect 148492 20412 148756 20422
rect 148548 20356 148596 20412
rect 148652 20356 148700 20412
rect 148492 20346 148756 20356
rect 148492 18844 148756 18854
rect 148548 18788 148596 18844
rect 148652 18788 148700 18844
rect 148492 18778 148756 18788
rect 148492 17276 148756 17286
rect 148548 17220 148596 17276
rect 148652 17220 148700 17276
rect 148492 17210 148756 17220
rect 148492 15708 148756 15718
rect 148548 15652 148596 15708
rect 148652 15652 148700 15708
rect 148492 15642 148756 15652
rect 148492 14140 148756 14150
rect 148548 14084 148596 14140
rect 148652 14084 148700 14140
rect 148492 14074 148756 14084
rect 148492 12572 148756 12582
rect 148548 12516 148596 12572
rect 148652 12516 148700 12572
rect 148492 12506 148756 12516
rect 148492 11004 148756 11014
rect 148548 10948 148596 11004
rect 148652 10948 148700 11004
rect 148492 10938 148756 10948
rect 148492 9436 148756 9446
rect 148548 9380 148596 9436
rect 148652 9380 148700 9436
rect 148492 9370 148756 9380
rect 148492 7868 148756 7878
rect 148548 7812 148596 7868
rect 148652 7812 148700 7868
rect 148492 7802 148756 7812
rect 148492 6300 148756 6310
rect 148548 6244 148596 6300
rect 148652 6244 148700 6300
rect 148492 6234 148756 6244
rect 148492 4732 148756 4742
rect 148548 4676 148596 4732
rect 148652 4676 148700 4732
rect 148492 4666 148756 4676
rect 147868 3266 147924 3276
rect 148492 3164 148756 3174
rect 148548 3108 148596 3164
rect 148652 3108 148700 3164
rect 148492 3098 148756 3108
rect 146076 2034 146132 2044
rect 145964 1138 146020 1148
rect 17276 700 17668 756
rect 18592 0 18704 800
rect 20272 0 20384 800
rect 21952 0 22064 800
rect 23632 0 23744 800
rect 25312 0 25424 800
rect 26992 0 27104 800
rect 28672 0 28784 800
rect 30352 0 30464 800
rect 32032 0 32144 800
rect 33712 0 33824 800
rect 35392 0 35504 800
rect 37072 0 37184 800
rect 38752 0 38864 800
rect 40432 0 40544 800
rect 42112 0 42224 800
rect 43792 0 43904 800
rect 45472 0 45584 800
rect 47152 0 47264 800
rect 48832 0 48944 800
rect 50512 0 50624 800
rect 52192 0 52304 800
rect 53872 0 53984 800
rect 55552 0 55664 800
rect 57232 0 57344 800
rect 58912 0 59024 800
rect 60592 0 60704 800
rect 62272 0 62384 800
rect 63952 0 64064 800
rect 65632 0 65744 800
rect 67312 0 67424 800
rect 68992 0 69104 800
rect 70672 0 70784 800
rect 72352 0 72464 800
rect 74032 0 74144 800
rect 75712 0 75824 800
rect 77392 0 77504 800
rect 79072 0 79184 800
rect 80752 0 80864 800
rect 82432 0 82544 800
rect 84112 0 84224 800
rect 85792 0 85904 800
rect 87472 0 87584 800
rect 89152 0 89264 800
rect 90832 0 90944 800
rect 92512 0 92624 800
rect 94192 0 94304 800
rect 95872 0 95984 800
rect 97552 0 97664 800
rect 99232 0 99344 800
rect 100912 0 101024 800
rect 102592 0 102704 800
rect 104272 0 104384 800
rect 105952 0 106064 800
rect 107632 0 107744 800
rect 109312 0 109424 800
rect 110992 0 111104 800
rect 112672 0 112784 800
rect 114352 0 114464 800
rect 116032 0 116144 800
rect 117712 0 117824 800
rect 119392 0 119504 800
rect 121072 0 121184 800
rect 122752 0 122864 800
rect 124432 0 124544 800
rect 126112 0 126224 800
rect 127792 0 127904 800
rect 129472 0 129584 800
rect 131152 0 131264 800
rect 132832 0 132944 800
rect 134512 0 134624 800
rect 136192 0 136304 800
rect 137872 0 137984 800
rect 139552 0 139664 800
rect 141232 0 141344 800
rect 142912 0 143024 800
rect 144592 0 144704 800
<< via2 >>
rect 147644 38780 147700 38836
rect 144508 37884 144564 37940
rect 19622 36874 19678 36876
rect 19622 36822 19624 36874
rect 19624 36822 19676 36874
rect 19676 36822 19678 36874
rect 19622 36820 19678 36822
rect 19726 36874 19782 36876
rect 19726 36822 19728 36874
rect 19728 36822 19780 36874
rect 19780 36822 19782 36874
rect 19726 36820 19782 36822
rect 19830 36874 19886 36876
rect 19830 36822 19832 36874
rect 19832 36822 19884 36874
rect 19884 36822 19886 36874
rect 19830 36820 19886 36822
rect 56442 36874 56498 36876
rect 56442 36822 56444 36874
rect 56444 36822 56496 36874
rect 56496 36822 56498 36874
rect 56442 36820 56498 36822
rect 56546 36874 56602 36876
rect 56546 36822 56548 36874
rect 56548 36822 56600 36874
rect 56600 36822 56602 36874
rect 56546 36820 56602 36822
rect 56650 36874 56706 36876
rect 56650 36822 56652 36874
rect 56652 36822 56704 36874
rect 56704 36822 56706 36874
rect 56650 36820 56706 36822
rect 93262 36874 93318 36876
rect 93262 36822 93264 36874
rect 93264 36822 93316 36874
rect 93316 36822 93318 36874
rect 93262 36820 93318 36822
rect 93366 36874 93422 36876
rect 93366 36822 93368 36874
rect 93368 36822 93420 36874
rect 93420 36822 93422 36874
rect 93366 36820 93422 36822
rect 93470 36874 93526 36876
rect 93470 36822 93472 36874
rect 93472 36822 93524 36874
rect 93524 36822 93526 36874
rect 93470 36820 93526 36822
rect 130082 36874 130138 36876
rect 130082 36822 130084 36874
rect 130084 36822 130136 36874
rect 130136 36822 130138 36874
rect 130082 36820 130138 36822
rect 130186 36874 130242 36876
rect 130186 36822 130188 36874
rect 130188 36822 130240 36874
rect 130240 36822 130242 36874
rect 130186 36820 130242 36822
rect 130290 36874 130346 36876
rect 130290 36822 130292 36874
rect 130292 36822 130344 36874
rect 130344 36822 130346 36874
rect 130290 36820 130346 36822
rect 139020 36204 139076 36260
rect 38032 36090 38088 36092
rect 38032 36038 38034 36090
rect 38034 36038 38086 36090
rect 38086 36038 38088 36090
rect 38032 36036 38088 36038
rect 38136 36090 38192 36092
rect 38136 36038 38138 36090
rect 38138 36038 38190 36090
rect 38190 36038 38192 36090
rect 38136 36036 38192 36038
rect 38240 36090 38296 36092
rect 38240 36038 38242 36090
rect 38242 36038 38294 36090
rect 38294 36038 38296 36090
rect 38240 36036 38296 36038
rect 74852 36090 74908 36092
rect 74852 36038 74854 36090
rect 74854 36038 74906 36090
rect 74906 36038 74908 36090
rect 74852 36036 74908 36038
rect 74956 36090 75012 36092
rect 74956 36038 74958 36090
rect 74958 36038 75010 36090
rect 75010 36038 75012 36090
rect 74956 36036 75012 36038
rect 75060 36090 75116 36092
rect 75060 36038 75062 36090
rect 75062 36038 75114 36090
rect 75114 36038 75116 36090
rect 75060 36036 75116 36038
rect 111672 36090 111728 36092
rect 111672 36038 111674 36090
rect 111674 36038 111726 36090
rect 111726 36038 111728 36090
rect 111672 36036 111728 36038
rect 111776 36090 111832 36092
rect 111776 36038 111778 36090
rect 111778 36038 111830 36090
rect 111830 36038 111832 36090
rect 111776 36036 111832 36038
rect 111880 36090 111936 36092
rect 111880 36038 111882 36090
rect 111882 36038 111934 36090
rect 111934 36038 111936 36090
rect 111880 36036 111936 36038
rect 19622 35306 19678 35308
rect 19622 35254 19624 35306
rect 19624 35254 19676 35306
rect 19676 35254 19678 35306
rect 19622 35252 19678 35254
rect 19726 35306 19782 35308
rect 19726 35254 19728 35306
rect 19728 35254 19780 35306
rect 19780 35254 19782 35306
rect 19726 35252 19782 35254
rect 19830 35306 19886 35308
rect 19830 35254 19832 35306
rect 19832 35254 19884 35306
rect 19884 35254 19886 35306
rect 19830 35252 19886 35254
rect 56442 35306 56498 35308
rect 56442 35254 56444 35306
rect 56444 35254 56496 35306
rect 56496 35254 56498 35306
rect 56442 35252 56498 35254
rect 56546 35306 56602 35308
rect 56546 35254 56548 35306
rect 56548 35254 56600 35306
rect 56600 35254 56602 35306
rect 56546 35252 56602 35254
rect 56650 35306 56706 35308
rect 56650 35254 56652 35306
rect 56652 35254 56704 35306
rect 56704 35254 56706 35306
rect 56650 35252 56706 35254
rect 93262 35306 93318 35308
rect 93262 35254 93264 35306
rect 93264 35254 93316 35306
rect 93316 35254 93318 35306
rect 93262 35252 93318 35254
rect 93366 35306 93422 35308
rect 93366 35254 93368 35306
rect 93368 35254 93420 35306
rect 93420 35254 93422 35306
rect 93366 35252 93422 35254
rect 93470 35306 93526 35308
rect 93470 35254 93472 35306
rect 93472 35254 93524 35306
rect 93524 35254 93526 35306
rect 93470 35252 93526 35254
rect 130082 35306 130138 35308
rect 130082 35254 130084 35306
rect 130084 35254 130136 35306
rect 130136 35254 130138 35306
rect 130082 35252 130138 35254
rect 130186 35306 130242 35308
rect 130186 35254 130188 35306
rect 130188 35254 130240 35306
rect 130240 35254 130242 35306
rect 130186 35252 130242 35254
rect 130290 35306 130346 35308
rect 130290 35254 130292 35306
rect 130292 35254 130344 35306
rect 130344 35254 130346 35306
rect 130290 35252 130346 35254
rect 38032 34522 38088 34524
rect 38032 34470 38034 34522
rect 38034 34470 38086 34522
rect 38086 34470 38088 34522
rect 38032 34468 38088 34470
rect 38136 34522 38192 34524
rect 38136 34470 38138 34522
rect 38138 34470 38190 34522
rect 38190 34470 38192 34522
rect 38136 34468 38192 34470
rect 38240 34522 38296 34524
rect 38240 34470 38242 34522
rect 38242 34470 38294 34522
rect 38294 34470 38296 34522
rect 38240 34468 38296 34470
rect 74852 34522 74908 34524
rect 74852 34470 74854 34522
rect 74854 34470 74906 34522
rect 74906 34470 74908 34522
rect 74852 34468 74908 34470
rect 74956 34522 75012 34524
rect 74956 34470 74958 34522
rect 74958 34470 75010 34522
rect 75010 34470 75012 34522
rect 74956 34468 75012 34470
rect 75060 34522 75116 34524
rect 75060 34470 75062 34522
rect 75062 34470 75114 34522
rect 75114 34470 75116 34522
rect 75060 34468 75116 34470
rect 111672 34522 111728 34524
rect 111672 34470 111674 34522
rect 111674 34470 111726 34522
rect 111726 34470 111728 34522
rect 111672 34468 111728 34470
rect 111776 34522 111832 34524
rect 111776 34470 111778 34522
rect 111778 34470 111830 34522
rect 111830 34470 111832 34522
rect 111776 34468 111832 34470
rect 111880 34522 111936 34524
rect 111880 34470 111882 34522
rect 111882 34470 111934 34522
rect 111934 34470 111936 34522
rect 111880 34468 111936 34470
rect 137340 33964 137396 34020
rect 19622 33738 19678 33740
rect 19622 33686 19624 33738
rect 19624 33686 19676 33738
rect 19676 33686 19678 33738
rect 19622 33684 19678 33686
rect 19726 33738 19782 33740
rect 19726 33686 19728 33738
rect 19728 33686 19780 33738
rect 19780 33686 19782 33738
rect 19726 33684 19782 33686
rect 19830 33738 19886 33740
rect 19830 33686 19832 33738
rect 19832 33686 19884 33738
rect 19884 33686 19886 33738
rect 19830 33684 19886 33686
rect 56442 33738 56498 33740
rect 56442 33686 56444 33738
rect 56444 33686 56496 33738
rect 56496 33686 56498 33738
rect 56442 33684 56498 33686
rect 56546 33738 56602 33740
rect 56546 33686 56548 33738
rect 56548 33686 56600 33738
rect 56600 33686 56602 33738
rect 56546 33684 56602 33686
rect 56650 33738 56706 33740
rect 56650 33686 56652 33738
rect 56652 33686 56704 33738
rect 56704 33686 56706 33738
rect 56650 33684 56706 33686
rect 93262 33738 93318 33740
rect 93262 33686 93264 33738
rect 93264 33686 93316 33738
rect 93316 33686 93318 33738
rect 93262 33684 93318 33686
rect 93366 33738 93422 33740
rect 93366 33686 93368 33738
rect 93368 33686 93420 33738
rect 93420 33686 93422 33738
rect 93366 33684 93422 33686
rect 93470 33738 93526 33740
rect 93470 33686 93472 33738
rect 93472 33686 93524 33738
rect 93524 33686 93526 33738
rect 93470 33684 93526 33686
rect 130082 33738 130138 33740
rect 130082 33686 130084 33738
rect 130084 33686 130136 33738
rect 130136 33686 130138 33738
rect 130082 33684 130138 33686
rect 130186 33738 130242 33740
rect 130186 33686 130188 33738
rect 130188 33686 130240 33738
rect 130240 33686 130242 33738
rect 130186 33684 130242 33686
rect 130290 33738 130346 33740
rect 130290 33686 130292 33738
rect 130292 33686 130344 33738
rect 130344 33686 130346 33738
rect 130290 33684 130346 33686
rect 134764 33068 134820 33124
rect 38032 32954 38088 32956
rect 38032 32902 38034 32954
rect 38034 32902 38086 32954
rect 38086 32902 38088 32954
rect 38032 32900 38088 32902
rect 38136 32954 38192 32956
rect 38136 32902 38138 32954
rect 38138 32902 38190 32954
rect 38190 32902 38192 32954
rect 38136 32900 38192 32902
rect 38240 32954 38296 32956
rect 38240 32902 38242 32954
rect 38242 32902 38294 32954
rect 38294 32902 38296 32954
rect 38240 32900 38296 32902
rect 74852 32954 74908 32956
rect 74852 32902 74854 32954
rect 74854 32902 74906 32954
rect 74906 32902 74908 32954
rect 74852 32900 74908 32902
rect 74956 32954 75012 32956
rect 74956 32902 74958 32954
rect 74958 32902 75010 32954
rect 75010 32902 75012 32954
rect 74956 32900 75012 32902
rect 75060 32954 75116 32956
rect 75060 32902 75062 32954
rect 75062 32902 75114 32954
rect 75114 32902 75116 32954
rect 75060 32900 75116 32902
rect 111672 32954 111728 32956
rect 111672 32902 111674 32954
rect 111674 32902 111726 32954
rect 111726 32902 111728 32954
rect 111672 32900 111728 32902
rect 111776 32954 111832 32956
rect 111776 32902 111778 32954
rect 111778 32902 111830 32954
rect 111830 32902 111832 32954
rect 111776 32900 111832 32902
rect 111880 32954 111936 32956
rect 111880 32902 111882 32954
rect 111882 32902 111934 32954
rect 111934 32902 111936 32954
rect 111880 32900 111936 32902
rect 19622 32170 19678 32172
rect 19622 32118 19624 32170
rect 19624 32118 19676 32170
rect 19676 32118 19678 32170
rect 19622 32116 19678 32118
rect 19726 32170 19782 32172
rect 19726 32118 19728 32170
rect 19728 32118 19780 32170
rect 19780 32118 19782 32170
rect 19726 32116 19782 32118
rect 19830 32170 19886 32172
rect 19830 32118 19832 32170
rect 19832 32118 19884 32170
rect 19884 32118 19886 32170
rect 19830 32116 19886 32118
rect 56442 32170 56498 32172
rect 56442 32118 56444 32170
rect 56444 32118 56496 32170
rect 56496 32118 56498 32170
rect 56442 32116 56498 32118
rect 56546 32170 56602 32172
rect 56546 32118 56548 32170
rect 56548 32118 56600 32170
rect 56600 32118 56602 32170
rect 56546 32116 56602 32118
rect 56650 32170 56706 32172
rect 56650 32118 56652 32170
rect 56652 32118 56704 32170
rect 56704 32118 56706 32170
rect 56650 32116 56706 32118
rect 93262 32170 93318 32172
rect 93262 32118 93264 32170
rect 93264 32118 93316 32170
rect 93316 32118 93318 32170
rect 93262 32116 93318 32118
rect 93366 32170 93422 32172
rect 93366 32118 93368 32170
rect 93368 32118 93420 32170
rect 93420 32118 93422 32170
rect 93366 32116 93422 32118
rect 93470 32170 93526 32172
rect 93470 32118 93472 32170
rect 93472 32118 93524 32170
rect 93524 32118 93526 32170
rect 93470 32116 93526 32118
rect 130082 32170 130138 32172
rect 130082 32118 130084 32170
rect 130084 32118 130136 32170
rect 130136 32118 130138 32170
rect 130082 32116 130138 32118
rect 130186 32170 130242 32172
rect 130186 32118 130188 32170
rect 130188 32118 130240 32170
rect 130240 32118 130242 32170
rect 130186 32116 130242 32118
rect 130290 32170 130346 32172
rect 130290 32118 130292 32170
rect 130292 32118 130344 32170
rect 130344 32118 130346 32170
rect 130290 32116 130346 32118
rect 133308 31500 133364 31556
rect 38032 31386 38088 31388
rect 38032 31334 38034 31386
rect 38034 31334 38086 31386
rect 38086 31334 38088 31386
rect 38032 31332 38088 31334
rect 38136 31386 38192 31388
rect 38136 31334 38138 31386
rect 38138 31334 38190 31386
rect 38190 31334 38192 31386
rect 38136 31332 38192 31334
rect 38240 31386 38296 31388
rect 38240 31334 38242 31386
rect 38242 31334 38294 31386
rect 38294 31334 38296 31386
rect 38240 31332 38296 31334
rect 74852 31386 74908 31388
rect 74852 31334 74854 31386
rect 74854 31334 74906 31386
rect 74906 31334 74908 31386
rect 74852 31332 74908 31334
rect 74956 31386 75012 31388
rect 74956 31334 74958 31386
rect 74958 31334 75010 31386
rect 75010 31334 75012 31386
rect 74956 31332 75012 31334
rect 75060 31386 75116 31388
rect 75060 31334 75062 31386
rect 75062 31334 75114 31386
rect 75114 31334 75116 31386
rect 75060 31332 75116 31334
rect 111672 31386 111728 31388
rect 111672 31334 111674 31386
rect 111674 31334 111726 31386
rect 111726 31334 111728 31386
rect 111672 31332 111728 31334
rect 111776 31386 111832 31388
rect 111776 31334 111778 31386
rect 111778 31334 111830 31386
rect 111830 31334 111832 31386
rect 111776 31332 111832 31334
rect 111880 31386 111936 31388
rect 111880 31334 111882 31386
rect 111882 31334 111934 31386
rect 111934 31334 111936 31386
rect 111880 31332 111936 31334
rect 131404 30828 131460 30884
rect 19622 30602 19678 30604
rect 19622 30550 19624 30602
rect 19624 30550 19676 30602
rect 19676 30550 19678 30602
rect 19622 30548 19678 30550
rect 19726 30602 19782 30604
rect 19726 30550 19728 30602
rect 19728 30550 19780 30602
rect 19780 30550 19782 30602
rect 19726 30548 19782 30550
rect 19830 30602 19886 30604
rect 19830 30550 19832 30602
rect 19832 30550 19884 30602
rect 19884 30550 19886 30602
rect 19830 30548 19886 30550
rect 56442 30602 56498 30604
rect 56442 30550 56444 30602
rect 56444 30550 56496 30602
rect 56496 30550 56498 30602
rect 56442 30548 56498 30550
rect 56546 30602 56602 30604
rect 56546 30550 56548 30602
rect 56548 30550 56600 30602
rect 56600 30550 56602 30602
rect 56546 30548 56602 30550
rect 56650 30602 56706 30604
rect 56650 30550 56652 30602
rect 56652 30550 56704 30602
rect 56704 30550 56706 30602
rect 56650 30548 56706 30550
rect 93262 30602 93318 30604
rect 93262 30550 93264 30602
rect 93264 30550 93316 30602
rect 93316 30550 93318 30602
rect 93262 30548 93318 30550
rect 93366 30602 93422 30604
rect 93366 30550 93368 30602
rect 93368 30550 93420 30602
rect 93420 30550 93422 30602
rect 93366 30548 93422 30550
rect 93470 30602 93526 30604
rect 93470 30550 93472 30602
rect 93472 30550 93524 30602
rect 93524 30550 93526 30602
rect 93470 30548 93526 30550
rect 130082 30602 130138 30604
rect 130082 30550 130084 30602
rect 130084 30550 130136 30602
rect 130136 30550 130138 30602
rect 130082 30548 130138 30550
rect 130186 30602 130242 30604
rect 130186 30550 130188 30602
rect 130188 30550 130240 30602
rect 130240 30550 130242 30602
rect 130186 30548 130242 30550
rect 130290 30602 130346 30604
rect 130290 30550 130292 30602
rect 130292 30550 130344 30602
rect 130344 30550 130346 30602
rect 130290 30548 130346 30550
rect 38032 29818 38088 29820
rect 38032 29766 38034 29818
rect 38034 29766 38086 29818
rect 38086 29766 38088 29818
rect 38032 29764 38088 29766
rect 38136 29818 38192 29820
rect 38136 29766 38138 29818
rect 38138 29766 38190 29818
rect 38190 29766 38192 29818
rect 38136 29764 38192 29766
rect 38240 29818 38296 29820
rect 38240 29766 38242 29818
rect 38242 29766 38294 29818
rect 38294 29766 38296 29818
rect 38240 29764 38296 29766
rect 74852 29818 74908 29820
rect 74852 29766 74854 29818
rect 74854 29766 74906 29818
rect 74906 29766 74908 29818
rect 74852 29764 74908 29766
rect 74956 29818 75012 29820
rect 74956 29766 74958 29818
rect 74958 29766 75010 29818
rect 75010 29766 75012 29818
rect 74956 29764 75012 29766
rect 75060 29818 75116 29820
rect 75060 29766 75062 29818
rect 75062 29766 75114 29818
rect 75114 29766 75116 29818
rect 75060 29764 75116 29766
rect 111672 29818 111728 29820
rect 111672 29766 111674 29818
rect 111674 29766 111726 29818
rect 111726 29766 111728 29818
rect 111672 29764 111728 29766
rect 111776 29818 111832 29820
rect 111776 29766 111778 29818
rect 111778 29766 111830 29818
rect 111830 29766 111832 29818
rect 111776 29764 111832 29766
rect 111880 29818 111936 29820
rect 111880 29766 111882 29818
rect 111882 29766 111934 29818
rect 111934 29766 111936 29818
rect 111880 29764 111936 29766
rect 127932 29260 127988 29316
rect 19622 29034 19678 29036
rect 19622 28982 19624 29034
rect 19624 28982 19676 29034
rect 19676 28982 19678 29034
rect 19622 28980 19678 28982
rect 19726 29034 19782 29036
rect 19726 28982 19728 29034
rect 19728 28982 19780 29034
rect 19780 28982 19782 29034
rect 19726 28980 19782 28982
rect 19830 29034 19886 29036
rect 19830 28982 19832 29034
rect 19832 28982 19884 29034
rect 19884 28982 19886 29034
rect 19830 28980 19886 28982
rect 56442 29034 56498 29036
rect 56442 28982 56444 29034
rect 56444 28982 56496 29034
rect 56496 28982 56498 29034
rect 56442 28980 56498 28982
rect 56546 29034 56602 29036
rect 56546 28982 56548 29034
rect 56548 28982 56600 29034
rect 56600 28982 56602 29034
rect 56546 28980 56602 28982
rect 56650 29034 56706 29036
rect 56650 28982 56652 29034
rect 56652 28982 56704 29034
rect 56704 28982 56706 29034
rect 56650 28980 56706 28982
rect 93262 29034 93318 29036
rect 93262 28982 93264 29034
rect 93264 28982 93316 29034
rect 93316 28982 93318 29034
rect 93262 28980 93318 28982
rect 93366 29034 93422 29036
rect 93366 28982 93368 29034
rect 93368 28982 93420 29034
rect 93420 28982 93422 29034
rect 93366 28980 93422 28982
rect 93470 29034 93526 29036
rect 93470 28982 93472 29034
rect 93472 28982 93524 29034
rect 93524 28982 93526 29034
rect 93470 28980 93526 28982
rect 38032 28250 38088 28252
rect 38032 28198 38034 28250
rect 38034 28198 38086 28250
rect 38086 28198 38088 28250
rect 38032 28196 38088 28198
rect 38136 28250 38192 28252
rect 38136 28198 38138 28250
rect 38138 28198 38190 28250
rect 38190 28198 38192 28250
rect 38136 28196 38192 28198
rect 38240 28250 38296 28252
rect 38240 28198 38242 28250
rect 38242 28198 38294 28250
rect 38294 28198 38296 28250
rect 38240 28196 38296 28198
rect 74852 28250 74908 28252
rect 74852 28198 74854 28250
rect 74854 28198 74906 28250
rect 74906 28198 74908 28250
rect 74852 28196 74908 28198
rect 74956 28250 75012 28252
rect 74956 28198 74958 28250
rect 74958 28198 75010 28250
rect 75010 28198 75012 28250
rect 74956 28196 75012 28198
rect 75060 28250 75116 28252
rect 75060 28198 75062 28250
rect 75062 28198 75114 28250
rect 75114 28198 75116 28250
rect 75060 28196 75116 28198
rect 111672 28250 111728 28252
rect 111672 28198 111674 28250
rect 111674 28198 111726 28250
rect 111726 28198 111728 28250
rect 111672 28196 111728 28198
rect 111776 28250 111832 28252
rect 111776 28198 111778 28250
rect 111778 28198 111830 28250
rect 111830 28198 111832 28250
rect 111776 28196 111832 28198
rect 111880 28250 111936 28252
rect 111880 28198 111882 28250
rect 111882 28198 111934 28250
rect 111934 28198 111936 28250
rect 111880 28196 111936 28198
rect 124908 27692 124964 27748
rect 19622 27466 19678 27468
rect 19622 27414 19624 27466
rect 19624 27414 19676 27466
rect 19676 27414 19678 27466
rect 19622 27412 19678 27414
rect 19726 27466 19782 27468
rect 19726 27414 19728 27466
rect 19728 27414 19780 27466
rect 19780 27414 19782 27466
rect 19726 27412 19782 27414
rect 19830 27466 19886 27468
rect 19830 27414 19832 27466
rect 19832 27414 19884 27466
rect 19884 27414 19886 27466
rect 19830 27412 19886 27414
rect 56442 27466 56498 27468
rect 56442 27414 56444 27466
rect 56444 27414 56496 27466
rect 56496 27414 56498 27466
rect 56442 27412 56498 27414
rect 56546 27466 56602 27468
rect 56546 27414 56548 27466
rect 56548 27414 56600 27466
rect 56600 27414 56602 27466
rect 56546 27412 56602 27414
rect 56650 27466 56706 27468
rect 56650 27414 56652 27466
rect 56652 27414 56704 27466
rect 56704 27414 56706 27466
rect 56650 27412 56706 27414
rect 93262 27466 93318 27468
rect 93262 27414 93264 27466
rect 93264 27414 93316 27466
rect 93316 27414 93318 27466
rect 93262 27412 93318 27414
rect 93366 27466 93422 27468
rect 93366 27414 93368 27466
rect 93368 27414 93420 27466
rect 93420 27414 93422 27466
rect 93366 27412 93422 27414
rect 93470 27466 93526 27468
rect 93470 27414 93472 27466
rect 93472 27414 93524 27466
rect 93524 27414 93526 27466
rect 93470 27412 93526 27414
rect 124124 26908 124180 26964
rect 38032 26682 38088 26684
rect 38032 26630 38034 26682
rect 38034 26630 38086 26682
rect 38086 26630 38088 26682
rect 38032 26628 38088 26630
rect 38136 26682 38192 26684
rect 38136 26630 38138 26682
rect 38138 26630 38190 26682
rect 38190 26630 38192 26682
rect 38136 26628 38192 26630
rect 38240 26682 38296 26684
rect 38240 26630 38242 26682
rect 38242 26630 38294 26682
rect 38294 26630 38296 26682
rect 38240 26628 38296 26630
rect 74852 26682 74908 26684
rect 74852 26630 74854 26682
rect 74854 26630 74906 26682
rect 74906 26630 74908 26682
rect 74852 26628 74908 26630
rect 74956 26682 75012 26684
rect 74956 26630 74958 26682
rect 74958 26630 75010 26682
rect 75010 26630 75012 26682
rect 74956 26628 75012 26630
rect 75060 26682 75116 26684
rect 75060 26630 75062 26682
rect 75062 26630 75114 26682
rect 75114 26630 75116 26682
rect 75060 26628 75116 26630
rect 111672 26682 111728 26684
rect 111672 26630 111674 26682
rect 111674 26630 111726 26682
rect 111726 26630 111728 26682
rect 111672 26628 111728 26630
rect 111776 26682 111832 26684
rect 111776 26630 111778 26682
rect 111778 26630 111830 26682
rect 111830 26630 111832 26682
rect 111776 26628 111832 26630
rect 111880 26682 111936 26684
rect 111880 26630 111882 26682
rect 111882 26630 111934 26682
rect 111934 26630 111936 26682
rect 111880 26628 111936 26630
rect 19622 25898 19678 25900
rect 19622 25846 19624 25898
rect 19624 25846 19676 25898
rect 19676 25846 19678 25898
rect 19622 25844 19678 25846
rect 19726 25898 19782 25900
rect 19726 25846 19728 25898
rect 19728 25846 19780 25898
rect 19780 25846 19782 25898
rect 19726 25844 19782 25846
rect 19830 25898 19886 25900
rect 19830 25846 19832 25898
rect 19832 25846 19884 25898
rect 19884 25846 19886 25898
rect 19830 25844 19886 25846
rect 56442 25898 56498 25900
rect 56442 25846 56444 25898
rect 56444 25846 56496 25898
rect 56496 25846 56498 25898
rect 56442 25844 56498 25846
rect 56546 25898 56602 25900
rect 56546 25846 56548 25898
rect 56548 25846 56600 25898
rect 56600 25846 56602 25898
rect 56546 25844 56602 25846
rect 56650 25898 56706 25900
rect 56650 25846 56652 25898
rect 56652 25846 56704 25898
rect 56704 25846 56706 25898
rect 56650 25844 56706 25846
rect 93262 25898 93318 25900
rect 93262 25846 93264 25898
rect 93264 25846 93316 25898
rect 93316 25846 93318 25898
rect 93262 25844 93318 25846
rect 93366 25898 93422 25900
rect 93366 25846 93368 25898
rect 93368 25846 93420 25898
rect 93420 25846 93422 25898
rect 93366 25844 93422 25846
rect 93470 25898 93526 25900
rect 93470 25846 93472 25898
rect 93472 25846 93524 25898
rect 93524 25846 93526 25898
rect 93470 25844 93526 25846
rect 38032 25114 38088 25116
rect 38032 25062 38034 25114
rect 38034 25062 38086 25114
rect 38086 25062 38088 25114
rect 38032 25060 38088 25062
rect 38136 25114 38192 25116
rect 38136 25062 38138 25114
rect 38138 25062 38190 25114
rect 38190 25062 38192 25114
rect 38136 25060 38192 25062
rect 38240 25114 38296 25116
rect 38240 25062 38242 25114
rect 38242 25062 38294 25114
rect 38294 25062 38296 25114
rect 38240 25060 38296 25062
rect 74852 25114 74908 25116
rect 74852 25062 74854 25114
rect 74854 25062 74906 25114
rect 74906 25062 74908 25114
rect 74852 25060 74908 25062
rect 74956 25114 75012 25116
rect 74956 25062 74958 25114
rect 74958 25062 75010 25114
rect 75010 25062 75012 25114
rect 74956 25060 75012 25062
rect 75060 25114 75116 25116
rect 75060 25062 75062 25114
rect 75062 25062 75114 25114
rect 75114 25062 75116 25114
rect 75060 25060 75116 25062
rect 111672 25114 111728 25116
rect 111672 25062 111674 25114
rect 111674 25062 111726 25114
rect 111726 25062 111728 25114
rect 111672 25060 111728 25062
rect 111776 25114 111832 25116
rect 111776 25062 111778 25114
rect 111778 25062 111830 25114
rect 111830 25062 111832 25114
rect 111776 25060 111832 25062
rect 111880 25114 111936 25116
rect 111880 25062 111882 25114
rect 111882 25062 111934 25114
rect 111934 25062 111936 25114
rect 111880 25060 111936 25062
rect 120092 25116 120148 25172
rect 119196 24556 119252 24612
rect 19622 24330 19678 24332
rect 19622 24278 19624 24330
rect 19624 24278 19676 24330
rect 19676 24278 19678 24330
rect 19622 24276 19678 24278
rect 19726 24330 19782 24332
rect 19726 24278 19728 24330
rect 19728 24278 19780 24330
rect 19780 24278 19782 24330
rect 19726 24276 19782 24278
rect 19830 24330 19886 24332
rect 19830 24278 19832 24330
rect 19832 24278 19884 24330
rect 19884 24278 19886 24330
rect 19830 24276 19886 24278
rect 56442 24330 56498 24332
rect 56442 24278 56444 24330
rect 56444 24278 56496 24330
rect 56496 24278 56498 24330
rect 56442 24276 56498 24278
rect 56546 24330 56602 24332
rect 56546 24278 56548 24330
rect 56548 24278 56600 24330
rect 56600 24278 56602 24330
rect 56546 24276 56602 24278
rect 56650 24330 56706 24332
rect 56650 24278 56652 24330
rect 56652 24278 56704 24330
rect 56704 24278 56706 24330
rect 56650 24276 56706 24278
rect 93262 24330 93318 24332
rect 93262 24278 93264 24330
rect 93264 24278 93316 24330
rect 93316 24278 93318 24330
rect 93262 24276 93318 24278
rect 93366 24330 93422 24332
rect 93366 24278 93368 24330
rect 93368 24278 93420 24330
rect 93420 24278 93422 24330
rect 93366 24276 93422 24278
rect 93470 24330 93526 24332
rect 93470 24278 93472 24330
rect 93472 24278 93524 24330
rect 93524 24278 93526 24330
rect 93470 24276 93526 24278
rect 38032 23546 38088 23548
rect 38032 23494 38034 23546
rect 38034 23494 38086 23546
rect 38086 23494 38088 23546
rect 38032 23492 38088 23494
rect 38136 23546 38192 23548
rect 38136 23494 38138 23546
rect 38138 23494 38190 23546
rect 38190 23494 38192 23546
rect 38136 23492 38192 23494
rect 38240 23546 38296 23548
rect 38240 23494 38242 23546
rect 38242 23494 38294 23546
rect 38294 23494 38296 23546
rect 38240 23492 38296 23494
rect 74852 23546 74908 23548
rect 74852 23494 74854 23546
rect 74854 23494 74906 23546
rect 74906 23494 74908 23546
rect 74852 23492 74908 23494
rect 74956 23546 75012 23548
rect 74956 23494 74958 23546
rect 74958 23494 75010 23546
rect 75010 23494 75012 23546
rect 74956 23492 75012 23494
rect 75060 23546 75116 23548
rect 75060 23494 75062 23546
rect 75062 23494 75114 23546
rect 75114 23494 75116 23546
rect 75060 23492 75116 23494
rect 111672 23546 111728 23548
rect 111672 23494 111674 23546
rect 111674 23494 111726 23546
rect 111726 23494 111728 23546
rect 111672 23492 111728 23494
rect 111776 23546 111832 23548
rect 111776 23494 111778 23546
rect 111778 23494 111830 23546
rect 111830 23494 111832 23546
rect 111776 23492 111832 23494
rect 111880 23546 111936 23548
rect 111880 23494 111882 23546
rect 111882 23494 111934 23546
rect 111934 23494 111936 23546
rect 111880 23492 111936 23494
rect 19622 22762 19678 22764
rect 19622 22710 19624 22762
rect 19624 22710 19676 22762
rect 19676 22710 19678 22762
rect 19622 22708 19678 22710
rect 19726 22762 19782 22764
rect 19726 22710 19728 22762
rect 19728 22710 19780 22762
rect 19780 22710 19782 22762
rect 19726 22708 19782 22710
rect 19830 22762 19886 22764
rect 19830 22710 19832 22762
rect 19832 22710 19884 22762
rect 19884 22710 19886 22762
rect 19830 22708 19886 22710
rect 56442 22762 56498 22764
rect 56442 22710 56444 22762
rect 56444 22710 56496 22762
rect 56496 22710 56498 22762
rect 56442 22708 56498 22710
rect 56546 22762 56602 22764
rect 56546 22710 56548 22762
rect 56548 22710 56600 22762
rect 56600 22710 56602 22762
rect 56546 22708 56602 22710
rect 56650 22762 56706 22764
rect 56650 22710 56652 22762
rect 56652 22710 56704 22762
rect 56704 22710 56706 22762
rect 56650 22708 56706 22710
rect 93262 22762 93318 22764
rect 93262 22710 93264 22762
rect 93264 22710 93316 22762
rect 93316 22710 93318 22762
rect 93262 22708 93318 22710
rect 93366 22762 93422 22764
rect 93366 22710 93368 22762
rect 93368 22710 93420 22762
rect 93420 22710 93422 22762
rect 93366 22708 93422 22710
rect 93470 22762 93526 22764
rect 93470 22710 93472 22762
rect 93472 22710 93524 22762
rect 93524 22710 93526 22762
rect 93470 22708 93526 22710
rect 113484 22092 113540 22148
rect 38032 21978 38088 21980
rect 38032 21926 38034 21978
rect 38034 21926 38086 21978
rect 38086 21926 38088 21978
rect 38032 21924 38088 21926
rect 38136 21978 38192 21980
rect 38136 21926 38138 21978
rect 38138 21926 38190 21978
rect 38190 21926 38192 21978
rect 38136 21924 38192 21926
rect 38240 21978 38296 21980
rect 38240 21926 38242 21978
rect 38242 21926 38294 21978
rect 38294 21926 38296 21978
rect 38240 21924 38296 21926
rect 74852 21978 74908 21980
rect 74852 21926 74854 21978
rect 74854 21926 74906 21978
rect 74906 21926 74908 21978
rect 74852 21924 74908 21926
rect 74956 21978 75012 21980
rect 74956 21926 74958 21978
rect 74958 21926 75010 21978
rect 75010 21926 75012 21978
rect 74956 21924 75012 21926
rect 75060 21978 75116 21980
rect 75060 21926 75062 21978
rect 75062 21926 75114 21978
rect 75114 21926 75116 21978
rect 75060 21924 75116 21926
rect 111672 21978 111728 21980
rect 111672 21926 111674 21978
rect 111674 21926 111726 21978
rect 111726 21926 111728 21978
rect 111672 21924 111728 21926
rect 111776 21978 111832 21980
rect 111776 21926 111778 21978
rect 111778 21926 111830 21978
rect 111830 21926 111832 21978
rect 111776 21924 111832 21926
rect 111880 21978 111936 21980
rect 111880 21926 111882 21978
rect 111882 21926 111934 21978
rect 111934 21926 111936 21978
rect 111880 21924 111936 21926
rect 19622 21194 19678 21196
rect 19622 21142 19624 21194
rect 19624 21142 19676 21194
rect 19676 21142 19678 21194
rect 19622 21140 19678 21142
rect 19726 21194 19782 21196
rect 19726 21142 19728 21194
rect 19728 21142 19780 21194
rect 19780 21142 19782 21194
rect 19726 21140 19782 21142
rect 19830 21194 19886 21196
rect 19830 21142 19832 21194
rect 19832 21142 19884 21194
rect 19884 21142 19886 21194
rect 19830 21140 19886 21142
rect 56442 21194 56498 21196
rect 56442 21142 56444 21194
rect 56444 21142 56496 21194
rect 56496 21142 56498 21194
rect 56442 21140 56498 21142
rect 56546 21194 56602 21196
rect 56546 21142 56548 21194
rect 56548 21142 56600 21194
rect 56600 21142 56602 21194
rect 56546 21140 56602 21142
rect 56650 21194 56706 21196
rect 56650 21142 56652 21194
rect 56652 21142 56704 21194
rect 56704 21142 56706 21194
rect 56650 21140 56706 21142
rect 93262 21194 93318 21196
rect 93262 21142 93264 21194
rect 93264 21142 93316 21194
rect 93316 21142 93318 21194
rect 93262 21140 93318 21142
rect 93366 21194 93422 21196
rect 93366 21142 93368 21194
rect 93368 21142 93420 21194
rect 93420 21142 93422 21194
rect 93366 21140 93422 21142
rect 93470 21194 93526 21196
rect 93470 21142 93472 21194
rect 93472 21142 93524 21194
rect 93524 21142 93526 21194
rect 93470 21140 93526 21142
rect 38032 20410 38088 20412
rect 38032 20358 38034 20410
rect 38034 20358 38086 20410
rect 38086 20358 38088 20410
rect 38032 20356 38088 20358
rect 38136 20410 38192 20412
rect 38136 20358 38138 20410
rect 38138 20358 38190 20410
rect 38190 20358 38192 20410
rect 38136 20356 38192 20358
rect 38240 20410 38296 20412
rect 38240 20358 38242 20410
rect 38242 20358 38294 20410
rect 38294 20358 38296 20410
rect 38240 20356 38296 20358
rect 74852 20410 74908 20412
rect 74852 20358 74854 20410
rect 74854 20358 74906 20410
rect 74906 20358 74908 20410
rect 74852 20356 74908 20358
rect 74956 20410 75012 20412
rect 74956 20358 74958 20410
rect 74958 20358 75010 20410
rect 75010 20358 75012 20410
rect 74956 20356 75012 20358
rect 75060 20410 75116 20412
rect 75060 20358 75062 20410
rect 75062 20358 75114 20410
rect 75114 20358 75116 20410
rect 75060 20356 75116 20358
rect 111672 20410 111728 20412
rect 111672 20358 111674 20410
rect 111674 20358 111726 20410
rect 111726 20358 111728 20410
rect 111672 20356 111728 20358
rect 111776 20410 111832 20412
rect 111776 20358 111778 20410
rect 111778 20358 111830 20410
rect 111830 20358 111832 20410
rect 111776 20356 111832 20358
rect 111880 20410 111936 20412
rect 111880 20358 111882 20410
rect 111882 20358 111934 20410
rect 111934 20358 111936 20410
rect 111880 20356 111936 20358
rect 19622 19626 19678 19628
rect 19622 19574 19624 19626
rect 19624 19574 19676 19626
rect 19676 19574 19678 19626
rect 19622 19572 19678 19574
rect 19726 19626 19782 19628
rect 19726 19574 19728 19626
rect 19728 19574 19780 19626
rect 19780 19574 19782 19626
rect 19726 19572 19782 19574
rect 19830 19626 19886 19628
rect 19830 19574 19832 19626
rect 19832 19574 19884 19626
rect 19884 19574 19886 19626
rect 19830 19572 19886 19574
rect 56442 19626 56498 19628
rect 56442 19574 56444 19626
rect 56444 19574 56496 19626
rect 56496 19574 56498 19626
rect 56442 19572 56498 19574
rect 56546 19626 56602 19628
rect 56546 19574 56548 19626
rect 56548 19574 56600 19626
rect 56600 19574 56602 19626
rect 56546 19572 56602 19574
rect 56650 19626 56706 19628
rect 56650 19574 56652 19626
rect 56652 19574 56704 19626
rect 56704 19574 56706 19626
rect 56650 19572 56706 19574
rect 93262 19626 93318 19628
rect 93262 19574 93264 19626
rect 93264 19574 93316 19626
rect 93316 19574 93318 19626
rect 93262 19572 93318 19574
rect 93366 19626 93422 19628
rect 93366 19574 93368 19626
rect 93368 19574 93420 19626
rect 93420 19574 93422 19626
rect 93366 19572 93422 19574
rect 93470 19626 93526 19628
rect 93470 19574 93472 19626
rect 93472 19574 93524 19626
rect 93524 19574 93526 19626
rect 93470 19572 93526 19574
rect 38032 18842 38088 18844
rect 38032 18790 38034 18842
rect 38034 18790 38086 18842
rect 38086 18790 38088 18842
rect 38032 18788 38088 18790
rect 38136 18842 38192 18844
rect 38136 18790 38138 18842
rect 38138 18790 38190 18842
rect 38190 18790 38192 18842
rect 38136 18788 38192 18790
rect 38240 18842 38296 18844
rect 38240 18790 38242 18842
rect 38242 18790 38294 18842
rect 38294 18790 38296 18842
rect 38240 18788 38296 18790
rect 74852 18842 74908 18844
rect 74852 18790 74854 18842
rect 74854 18790 74906 18842
rect 74906 18790 74908 18842
rect 74852 18788 74908 18790
rect 74956 18842 75012 18844
rect 74956 18790 74958 18842
rect 74958 18790 75010 18842
rect 75010 18790 75012 18842
rect 74956 18788 75012 18790
rect 75060 18842 75116 18844
rect 75060 18790 75062 18842
rect 75062 18790 75114 18842
rect 75114 18790 75116 18842
rect 75060 18788 75116 18790
rect 111672 18842 111728 18844
rect 111672 18790 111674 18842
rect 111674 18790 111726 18842
rect 111726 18790 111728 18842
rect 111672 18788 111728 18790
rect 111776 18842 111832 18844
rect 111776 18790 111778 18842
rect 111778 18790 111830 18842
rect 111830 18790 111832 18842
rect 111776 18788 111832 18790
rect 111880 18842 111936 18844
rect 111880 18790 111882 18842
rect 111882 18790 111934 18842
rect 111934 18790 111936 18842
rect 111880 18788 111936 18790
rect 111580 18674 111636 18676
rect 111580 18622 111582 18674
rect 111582 18622 111634 18674
rect 111634 18622 111636 18674
rect 111580 18620 111636 18622
rect 19622 18058 19678 18060
rect 19622 18006 19624 18058
rect 19624 18006 19676 18058
rect 19676 18006 19678 18058
rect 19622 18004 19678 18006
rect 19726 18058 19782 18060
rect 19726 18006 19728 18058
rect 19728 18006 19780 18058
rect 19780 18006 19782 18058
rect 19726 18004 19782 18006
rect 19830 18058 19886 18060
rect 19830 18006 19832 18058
rect 19832 18006 19884 18058
rect 19884 18006 19886 18058
rect 19830 18004 19886 18006
rect 56442 18058 56498 18060
rect 56442 18006 56444 18058
rect 56444 18006 56496 18058
rect 56496 18006 56498 18058
rect 56442 18004 56498 18006
rect 56546 18058 56602 18060
rect 56546 18006 56548 18058
rect 56548 18006 56600 18058
rect 56600 18006 56602 18058
rect 56546 18004 56602 18006
rect 56650 18058 56706 18060
rect 56650 18006 56652 18058
rect 56652 18006 56704 18058
rect 56704 18006 56706 18058
rect 56650 18004 56706 18006
rect 93262 18058 93318 18060
rect 93262 18006 93264 18058
rect 93264 18006 93316 18058
rect 93316 18006 93318 18058
rect 93262 18004 93318 18006
rect 93366 18058 93422 18060
rect 93366 18006 93368 18058
rect 93368 18006 93420 18058
rect 93420 18006 93422 18058
rect 93366 18004 93422 18006
rect 93470 18058 93526 18060
rect 93470 18006 93472 18058
rect 93472 18006 93524 18058
rect 93524 18006 93526 18058
rect 93470 18004 93526 18006
rect 106652 17388 106708 17444
rect 38032 17274 38088 17276
rect 38032 17222 38034 17274
rect 38034 17222 38086 17274
rect 38086 17222 38088 17274
rect 38032 17220 38088 17222
rect 38136 17274 38192 17276
rect 38136 17222 38138 17274
rect 38138 17222 38190 17274
rect 38190 17222 38192 17274
rect 38136 17220 38192 17222
rect 38240 17274 38296 17276
rect 38240 17222 38242 17274
rect 38242 17222 38294 17274
rect 38294 17222 38296 17274
rect 38240 17220 38296 17222
rect 74852 17274 74908 17276
rect 74852 17222 74854 17274
rect 74854 17222 74906 17274
rect 74906 17222 74908 17274
rect 74852 17220 74908 17222
rect 74956 17274 75012 17276
rect 74956 17222 74958 17274
rect 74958 17222 75010 17274
rect 75010 17222 75012 17274
rect 74956 17220 75012 17222
rect 75060 17274 75116 17276
rect 75060 17222 75062 17274
rect 75062 17222 75114 17274
rect 75114 17222 75116 17274
rect 75060 17220 75116 17222
rect 104524 16828 104580 16884
rect 19622 16490 19678 16492
rect 19622 16438 19624 16490
rect 19624 16438 19676 16490
rect 19676 16438 19678 16490
rect 19622 16436 19678 16438
rect 19726 16490 19782 16492
rect 19726 16438 19728 16490
rect 19728 16438 19780 16490
rect 19780 16438 19782 16490
rect 19726 16436 19782 16438
rect 19830 16490 19886 16492
rect 19830 16438 19832 16490
rect 19832 16438 19884 16490
rect 19884 16438 19886 16490
rect 19830 16436 19886 16438
rect 56442 16490 56498 16492
rect 56442 16438 56444 16490
rect 56444 16438 56496 16490
rect 56496 16438 56498 16490
rect 56442 16436 56498 16438
rect 56546 16490 56602 16492
rect 56546 16438 56548 16490
rect 56548 16438 56600 16490
rect 56600 16438 56602 16490
rect 56546 16436 56602 16438
rect 56650 16490 56706 16492
rect 56650 16438 56652 16490
rect 56652 16438 56704 16490
rect 56704 16438 56706 16490
rect 56650 16436 56706 16438
rect 93262 16490 93318 16492
rect 93262 16438 93264 16490
rect 93264 16438 93316 16490
rect 93316 16438 93318 16490
rect 93262 16436 93318 16438
rect 93366 16490 93422 16492
rect 93366 16438 93368 16490
rect 93368 16438 93420 16490
rect 93420 16438 93422 16490
rect 93366 16436 93422 16438
rect 93470 16490 93526 16492
rect 93470 16438 93472 16490
rect 93472 16438 93524 16490
rect 93524 16438 93526 16490
rect 93470 16436 93526 16438
rect 103628 15820 103684 15876
rect 38032 15706 38088 15708
rect 38032 15654 38034 15706
rect 38034 15654 38086 15706
rect 38086 15654 38088 15706
rect 38032 15652 38088 15654
rect 38136 15706 38192 15708
rect 38136 15654 38138 15706
rect 38138 15654 38190 15706
rect 38190 15654 38192 15706
rect 38136 15652 38192 15654
rect 38240 15706 38296 15708
rect 38240 15654 38242 15706
rect 38242 15654 38294 15706
rect 38294 15654 38296 15706
rect 38240 15652 38296 15654
rect 74852 15706 74908 15708
rect 74852 15654 74854 15706
rect 74854 15654 74906 15706
rect 74906 15654 74908 15706
rect 74852 15652 74908 15654
rect 74956 15706 75012 15708
rect 74956 15654 74958 15706
rect 74958 15654 75010 15706
rect 75010 15654 75012 15706
rect 74956 15652 75012 15654
rect 75060 15706 75116 15708
rect 75060 15654 75062 15706
rect 75062 15654 75114 15706
rect 75114 15654 75116 15706
rect 75060 15652 75116 15654
rect 19622 14922 19678 14924
rect 19622 14870 19624 14922
rect 19624 14870 19676 14922
rect 19676 14870 19678 14922
rect 19622 14868 19678 14870
rect 19726 14922 19782 14924
rect 19726 14870 19728 14922
rect 19728 14870 19780 14922
rect 19780 14870 19782 14922
rect 19726 14868 19782 14870
rect 19830 14922 19886 14924
rect 19830 14870 19832 14922
rect 19832 14870 19884 14922
rect 19884 14870 19886 14922
rect 19830 14868 19886 14870
rect 56442 14922 56498 14924
rect 56442 14870 56444 14922
rect 56444 14870 56496 14922
rect 56496 14870 56498 14922
rect 56442 14868 56498 14870
rect 56546 14922 56602 14924
rect 56546 14870 56548 14922
rect 56548 14870 56600 14922
rect 56600 14870 56602 14922
rect 56546 14868 56602 14870
rect 56650 14922 56706 14924
rect 56650 14870 56652 14922
rect 56652 14870 56704 14922
rect 56704 14870 56706 14922
rect 56650 14868 56706 14870
rect 93262 14922 93318 14924
rect 93262 14870 93264 14922
rect 93264 14870 93316 14922
rect 93316 14870 93318 14922
rect 93262 14868 93318 14870
rect 93366 14922 93422 14924
rect 93366 14870 93368 14922
rect 93368 14870 93420 14922
rect 93420 14870 93422 14922
rect 93366 14868 93422 14870
rect 93470 14922 93526 14924
rect 93470 14870 93472 14922
rect 93472 14870 93524 14922
rect 93524 14870 93526 14922
rect 93470 14868 93526 14870
rect 100492 14252 100548 14308
rect 38032 14138 38088 14140
rect 38032 14086 38034 14138
rect 38034 14086 38086 14138
rect 38086 14086 38088 14138
rect 38032 14084 38088 14086
rect 38136 14138 38192 14140
rect 38136 14086 38138 14138
rect 38138 14086 38190 14138
rect 38190 14086 38192 14138
rect 38136 14084 38192 14086
rect 38240 14138 38296 14140
rect 38240 14086 38242 14138
rect 38242 14086 38294 14138
rect 38294 14086 38296 14138
rect 38240 14084 38296 14086
rect 74852 14138 74908 14140
rect 74852 14086 74854 14138
rect 74854 14086 74906 14138
rect 74906 14086 74908 14138
rect 74852 14084 74908 14086
rect 74956 14138 75012 14140
rect 74956 14086 74958 14138
rect 74958 14086 75010 14138
rect 75010 14086 75012 14138
rect 74956 14084 75012 14086
rect 75060 14138 75116 14140
rect 75060 14086 75062 14138
rect 75062 14086 75114 14138
rect 75114 14086 75116 14138
rect 75060 14084 75116 14086
rect 19622 13354 19678 13356
rect 19622 13302 19624 13354
rect 19624 13302 19676 13354
rect 19676 13302 19678 13354
rect 19622 13300 19678 13302
rect 19726 13354 19782 13356
rect 19726 13302 19728 13354
rect 19728 13302 19780 13354
rect 19780 13302 19782 13354
rect 19726 13300 19782 13302
rect 19830 13354 19886 13356
rect 19830 13302 19832 13354
rect 19832 13302 19884 13354
rect 19884 13302 19886 13354
rect 19830 13300 19886 13302
rect 56442 13354 56498 13356
rect 56442 13302 56444 13354
rect 56444 13302 56496 13354
rect 56496 13302 56498 13354
rect 56442 13300 56498 13302
rect 56546 13354 56602 13356
rect 56546 13302 56548 13354
rect 56548 13302 56600 13354
rect 56600 13302 56602 13354
rect 56546 13300 56602 13302
rect 56650 13354 56706 13356
rect 56650 13302 56652 13354
rect 56652 13302 56704 13354
rect 56704 13302 56706 13354
rect 56650 13300 56706 13302
rect 93262 13354 93318 13356
rect 93262 13302 93264 13354
rect 93264 13302 93316 13354
rect 93316 13302 93318 13354
rect 93262 13300 93318 13302
rect 93366 13354 93422 13356
rect 93366 13302 93368 13354
rect 93368 13302 93420 13354
rect 93420 13302 93422 13354
rect 93366 13300 93422 13302
rect 93470 13354 93526 13356
rect 93470 13302 93472 13354
rect 93472 13302 93524 13354
rect 93524 13302 93526 13354
rect 93470 13300 93526 13302
rect 100044 12796 100100 12852
rect 38032 12570 38088 12572
rect 38032 12518 38034 12570
rect 38034 12518 38086 12570
rect 38086 12518 38088 12570
rect 38032 12516 38088 12518
rect 38136 12570 38192 12572
rect 38136 12518 38138 12570
rect 38138 12518 38190 12570
rect 38190 12518 38192 12570
rect 38136 12516 38192 12518
rect 38240 12570 38296 12572
rect 38240 12518 38242 12570
rect 38242 12518 38294 12570
rect 38294 12518 38296 12570
rect 38240 12516 38296 12518
rect 74852 12570 74908 12572
rect 74852 12518 74854 12570
rect 74854 12518 74906 12570
rect 74906 12518 74908 12570
rect 74852 12516 74908 12518
rect 74956 12570 75012 12572
rect 74956 12518 74958 12570
rect 74958 12518 75010 12570
rect 75010 12518 75012 12570
rect 74956 12516 75012 12518
rect 75060 12570 75116 12572
rect 75060 12518 75062 12570
rect 75062 12518 75114 12570
rect 75114 12518 75116 12570
rect 75060 12516 75116 12518
rect 71372 12348 71428 12404
rect 63868 11900 63924 11956
rect 19622 11786 19678 11788
rect 19622 11734 19624 11786
rect 19624 11734 19676 11786
rect 19676 11734 19678 11786
rect 19622 11732 19678 11734
rect 19726 11786 19782 11788
rect 19726 11734 19728 11786
rect 19728 11734 19780 11786
rect 19780 11734 19782 11786
rect 19726 11732 19782 11734
rect 19830 11786 19886 11788
rect 19830 11734 19832 11786
rect 19832 11734 19884 11786
rect 19884 11734 19886 11786
rect 19830 11732 19886 11734
rect 56442 11786 56498 11788
rect 56442 11734 56444 11786
rect 56444 11734 56496 11786
rect 56496 11734 56498 11786
rect 56442 11732 56498 11734
rect 56546 11786 56602 11788
rect 56546 11734 56548 11786
rect 56548 11734 56600 11786
rect 56600 11734 56602 11786
rect 56546 11732 56602 11734
rect 56650 11786 56706 11788
rect 56650 11734 56652 11786
rect 56652 11734 56704 11786
rect 56704 11734 56706 11786
rect 56650 11732 56706 11734
rect 38032 11002 38088 11004
rect 38032 10950 38034 11002
rect 38034 10950 38086 11002
rect 38086 10950 38088 11002
rect 38032 10948 38088 10950
rect 38136 11002 38192 11004
rect 38136 10950 38138 11002
rect 38138 10950 38190 11002
rect 38190 10950 38192 11002
rect 38136 10948 38192 10950
rect 38240 11002 38296 11004
rect 38240 10950 38242 11002
rect 38242 10950 38294 11002
rect 38294 10950 38296 11002
rect 38240 10948 38296 10950
rect 53900 10668 53956 10724
rect 32396 10556 32452 10612
rect 17052 10332 17108 10388
rect 12124 8988 12180 9044
rect 10780 7308 10836 7364
rect 9996 5068 10052 5124
rect 8764 4508 8820 4564
rect 8316 4338 8372 4340
rect 8316 4286 8318 4338
rect 8318 4286 8370 4338
rect 8370 4286 8372 4338
rect 8316 4284 8372 4286
rect 5180 3388 5236 3444
rect 5852 3442 5908 3444
rect 5852 3390 5854 3442
rect 5854 3390 5906 3442
rect 5906 3390 5908 3442
rect 5852 3388 5908 3390
rect 6972 3276 7028 3332
rect 9772 4562 9828 4564
rect 9772 4510 9774 4562
rect 9774 4510 9826 4562
rect 9826 4510 9828 4562
rect 9772 4508 9828 4510
rect 8876 4338 8932 4340
rect 8876 4286 8878 4338
rect 8878 4286 8930 4338
rect 8930 4286 8932 4338
rect 8876 4284 8932 4286
rect 10780 4508 10836 4564
rect 11004 4508 11060 4564
rect 9996 4284 10052 4340
rect 11340 4562 11396 4564
rect 11340 4510 11342 4562
rect 11342 4510 11394 4562
rect 11394 4510 11396 4562
rect 11340 4508 11396 4510
rect 15036 8876 15092 8932
rect 12124 4508 12180 4564
rect 13020 4562 13076 4564
rect 13020 4510 13022 4562
rect 13022 4510 13074 4562
rect 13074 4510 13076 4562
rect 13020 4508 13076 4510
rect 15036 4508 15092 4564
rect 19622 10218 19678 10220
rect 19622 10166 19624 10218
rect 19624 10166 19676 10218
rect 19676 10166 19678 10218
rect 19622 10164 19678 10166
rect 19726 10218 19782 10220
rect 19726 10166 19728 10218
rect 19728 10166 19780 10218
rect 19780 10166 19782 10218
rect 19726 10164 19782 10166
rect 19830 10218 19886 10220
rect 19830 10166 19832 10218
rect 19832 10166 19884 10218
rect 19884 10166 19886 10218
rect 19830 10164 19886 10166
rect 19622 8650 19678 8652
rect 19622 8598 19624 8650
rect 19624 8598 19676 8650
rect 19676 8598 19678 8650
rect 19622 8596 19678 8598
rect 19726 8650 19782 8652
rect 19726 8598 19728 8650
rect 19728 8598 19780 8650
rect 19780 8598 19782 8650
rect 19726 8596 19782 8598
rect 19830 8650 19886 8652
rect 19830 8598 19832 8650
rect 19832 8598 19884 8650
rect 19884 8598 19886 8650
rect 19830 8596 19886 8598
rect 19622 7082 19678 7084
rect 19622 7030 19624 7082
rect 19624 7030 19676 7082
rect 19676 7030 19678 7082
rect 19622 7028 19678 7030
rect 19726 7082 19782 7084
rect 19726 7030 19728 7082
rect 19728 7030 19780 7082
rect 19780 7030 19782 7082
rect 19726 7028 19782 7030
rect 19830 7082 19886 7084
rect 19830 7030 19832 7082
rect 19832 7030 19884 7082
rect 19884 7030 19886 7082
rect 19830 7028 19886 7030
rect 30044 5852 30100 5908
rect 28588 5628 28644 5684
rect 19622 5514 19678 5516
rect 19622 5462 19624 5514
rect 19624 5462 19676 5514
rect 19676 5462 19678 5514
rect 19622 5460 19678 5462
rect 19726 5514 19782 5516
rect 19726 5462 19728 5514
rect 19728 5462 19780 5514
rect 19780 5462 19782 5514
rect 19726 5460 19782 5462
rect 19830 5514 19886 5516
rect 19830 5462 19832 5514
rect 19832 5462 19884 5514
rect 19884 5462 19886 5514
rect 19830 5460 19886 5462
rect 14924 3724 14980 3780
rect 15148 3724 15204 3780
rect 27132 5292 27188 5348
rect 18284 3612 18340 3668
rect 20076 4060 20132 4116
rect 20524 4060 20580 4116
rect 19622 3946 19678 3948
rect 19622 3894 19624 3946
rect 19624 3894 19676 3946
rect 19676 3894 19678 3946
rect 19622 3892 19678 3894
rect 19726 3946 19782 3948
rect 19726 3894 19728 3946
rect 19728 3894 19780 3946
rect 19780 3894 19782 3946
rect 19726 3892 19782 3894
rect 19830 3946 19886 3948
rect 19830 3894 19832 3946
rect 19832 3894 19884 3946
rect 19884 3894 19886 3946
rect 19830 3892 19886 3894
rect 20636 3836 20692 3892
rect 18732 3612 18788 3668
rect 21420 3836 21476 3892
rect 23660 3388 23716 3444
rect 23772 2380 23828 2436
rect 25228 3442 25284 3444
rect 25228 3390 25230 3442
rect 25230 3390 25282 3442
rect 25282 3390 25284 3442
rect 25228 3388 25284 3390
rect 24556 1596 24612 1652
rect 28700 3500 28756 3556
rect 27132 3442 27188 3444
rect 27132 3390 27134 3442
rect 27134 3390 27186 3442
rect 27186 3390 27188 3442
rect 27132 3388 27188 3390
rect 30268 3554 30324 3556
rect 30268 3502 30270 3554
rect 30270 3502 30322 3554
rect 30322 3502 30324 3554
rect 30268 3500 30324 3502
rect 29148 3442 29204 3444
rect 29148 3390 29150 3442
rect 29150 3390 29202 3442
rect 29202 3390 29204 3442
rect 29148 3388 29204 3390
rect 31388 3442 31444 3444
rect 31388 3390 31390 3442
rect 31390 3390 31442 3442
rect 31442 3390 31444 3442
rect 31388 3388 31444 3390
rect 38032 9434 38088 9436
rect 38032 9382 38034 9434
rect 38034 9382 38086 9434
rect 38086 9382 38088 9434
rect 38032 9380 38088 9382
rect 38136 9434 38192 9436
rect 38136 9382 38138 9434
rect 38138 9382 38190 9434
rect 38190 9382 38192 9434
rect 38136 9380 38192 9382
rect 38240 9434 38296 9436
rect 38240 9382 38242 9434
rect 38242 9382 38294 9434
rect 38294 9382 38296 9434
rect 38240 9380 38296 9382
rect 47180 9100 47236 9156
rect 38032 7866 38088 7868
rect 38032 7814 38034 7866
rect 38034 7814 38086 7866
rect 38086 7814 38088 7866
rect 38032 7812 38088 7814
rect 38136 7866 38192 7868
rect 38136 7814 38138 7866
rect 38138 7814 38190 7866
rect 38190 7814 38192 7866
rect 38136 7812 38192 7814
rect 38240 7866 38296 7868
rect 38240 7814 38242 7866
rect 38242 7814 38294 7866
rect 38294 7814 38296 7866
rect 38240 7812 38296 7814
rect 36316 7196 36372 7252
rect 32956 4226 33012 4228
rect 32956 4174 32958 4226
rect 32958 4174 33010 4226
rect 33010 4174 33012 4226
rect 32956 4172 33012 4174
rect 33740 4172 33796 4228
rect 31948 2268 32004 2324
rect 32060 3388 32116 3444
rect 33068 3442 33124 3444
rect 33068 3390 33070 3442
rect 33070 3390 33122 3442
rect 33122 3390 33124 3442
rect 33068 3388 33124 3390
rect 35420 3388 35476 3444
rect 40348 6748 40404 6804
rect 38032 6298 38088 6300
rect 38032 6246 38034 6298
rect 38034 6246 38086 6298
rect 38086 6246 38088 6298
rect 38032 6244 38088 6246
rect 38136 6298 38192 6300
rect 38136 6246 38138 6298
rect 38138 6246 38190 6298
rect 38190 6246 38192 6298
rect 38136 6244 38192 6246
rect 38240 6298 38296 6300
rect 38240 6246 38242 6298
rect 38242 6246 38294 6298
rect 38294 6246 38296 6298
rect 38240 6244 38296 6246
rect 38032 4730 38088 4732
rect 38032 4678 38034 4730
rect 38034 4678 38086 4730
rect 38086 4678 38088 4730
rect 38032 4676 38088 4678
rect 38136 4730 38192 4732
rect 38136 4678 38138 4730
rect 38138 4678 38190 4730
rect 38190 4678 38192 4730
rect 38136 4676 38192 4678
rect 38240 4730 38296 4732
rect 38240 4678 38242 4730
rect 38242 4678 38294 4730
rect 38294 4678 38296 4730
rect 38240 4676 38296 4678
rect 36988 3442 37044 3444
rect 36988 3390 36990 3442
rect 36990 3390 37042 3442
rect 37042 3390 37044 3442
rect 36988 3388 37044 3390
rect 35644 812 35700 868
rect 38032 3162 38088 3164
rect 38032 3110 38034 3162
rect 38034 3110 38086 3162
rect 38086 3110 38088 3162
rect 38032 3108 38088 3110
rect 38136 3162 38192 3164
rect 38136 3110 38138 3162
rect 38138 3110 38190 3162
rect 38190 3110 38192 3162
rect 38136 3108 38192 3110
rect 38240 3162 38296 3164
rect 38240 3110 38242 3162
rect 38242 3110 38294 3162
rect 38294 3110 38296 3162
rect 38240 3108 38296 3110
rect 40796 4396 40852 4452
rect 41692 4450 41748 4452
rect 41692 4398 41694 4450
rect 41694 4398 41746 4450
rect 41746 4398 41748 4450
rect 41692 4396 41748 4398
rect 38668 2604 38724 2660
rect 38892 3442 38948 3444
rect 38892 3390 38894 3442
rect 38894 3390 38946 3442
rect 38946 3390 38948 3442
rect 38892 3388 38948 3390
rect 40908 3442 40964 3444
rect 40908 3390 40910 3442
rect 40910 3390 40962 3442
rect 40962 3390 40964 3442
rect 40908 3388 40964 3390
rect 43036 2828 43092 2884
rect 43708 1036 43764 1092
rect 43820 3388 43876 3444
rect 45388 3442 45444 3444
rect 45388 3390 45390 3442
rect 45390 3390 45442 3442
rect 45442 3390 45444 3442
rect 45388 3388 45444 3390
rect 45164 1484 45220 1540
rect 50988 7532 51044 7588
rect 48860 4396 48916 4452
rect 49644 4450 49700 4452
rect 49644 4398 49646 4450
rect 49646 4398 49698 4450
rect 49698 4398 49700 4450
rect 49644 4396 49700 4398
rect 47180 3388 47236 3444
rect 48748 3442 48804 3444
rect 48748 3390 48750 3442
rect 48750 3390 48802 3442
rect 48802 3390 48804 3442
rect 48748 3388 48804 3390
rect 48076 2716 48132 2772
rect 50652 3442 50708 3444
rect 50652 3390 50654 3442
rect 50654 3390 50706 3442
rect 50706 3390 50708 3442
rect 50652 3388 50708 3390
rect 52108 1260 52164 1316
rect 56442 10218 56498 10220
rect 56442 10166 56444 10218
rect 56444 10166 56496 10218
rect 56496 10166 56498 10218
rect 56442 10164 56498 10166
rect 56546 10218 56602 10220
rect 56546 10166 56548 10218
rect 56548 10166 56600 10218
rect 56600 10166 56602 10218
rect 56546 10164 56602 10166
rect 56650 10218 56706 10220
rect 56650 10166 56652 10218
rect 56652 10166 56704 10218
rect 56704 10166 56706 10218
rect 56650 10164 56706 10166
rect 56442 8650 56498 8652
rect 56442 8598 56444 8650
rect 56444 8598 56496 8650
rect 56496 8598 56498 8650
rect 56442 8596 56498 8598
rect 56546 8650 56602 8652
rect 56546 8598 56548 8650
rect 56548 8598 56600 8650
rect 56600 8598 56602 8650
rect 56546 8596 56602 8598
rect 56650 8650 56706 8652
rect 56650 8598 56652 8650
rect 56652 8598 56704 8650
rect 56704 8598 56706 8650
rect 56650 8596 56706 8598
rect 57036 8428 57092 8484
rect 56442 7082 56498 7084
rect 56442 7030 56444 7082
rect 56444 7030 56496 7082
rect 56496 7030 56498 7082
rect 56442 7028 56498 7030
rect 56546 7082 56602 7084
rect 56546 7030 56548 7082
rect 56548 7030 56600 7082
rect 56600 7030 56602 7082
rect 56546 7028 56602 7030
rect 56650 7082 56706 7084
rect 56650 7030 56652 7082
rect 56652 7030 56704 7082
rect 56704 7030 56706 7082
rect 56650 7028 56706 7030
rect 56442 5514 56498 5516
rect 56442 5462 56444 5514
rect 56444 5462 56496 5514
rect 56496 5462 56498 5514
rect 56442 5460 56498 5462
rect 56546 5514 56602 5516
rect 56546 5462 56548 5514
rect 56548 5462 56600 5514
rect 56600 5462 56602 5514
rect 56546 5460 56602 5462
rect 56650 5514 56706 5516
rect 56650 5462 56652 5514
rect 56652 5462 56704 5514
rect 56704 5462 56706 5514
rect 56650 5460 56706 5462
rect 52668 3442 52724 3444
rect 52668 3390 52670 3442
rect 52670 3390 52722 3442
rect 52722 3390 52724 3442
rect 52668 3388 52724 3390
rect 55468 2940 55524 2996
rect 59836 6860 59892 6916
rect 56442 3946 56498 3948
rect 56442 3894 56444 3946
rect 56444 3894 56496 3946
rect 56496 3894 56498 3946
rect 56442 3892 56498 3894
rect 56546 3946 56602 3948
rect 56546 3894 56548 3946
rect 56548 3894 56600 3946
rect 56600 3894 56602 3946
rect 56546 3892 56602 3894
rect 56650 3946 56706 3948
rect 56650 3894 56652 3946
rect 56652 3894 56704 3946
rect 56704 3894 56706 3946
rect 56650 3892 56706 3894
rect 58940 3388 58996 3444
rect 63756 4844 63812 4900
rect 60508 3442 60564 3444
rect 60508 3390 60510 3442
rect 60510 3390 60562 3442
rect 60562 3390 60564 3442
rect 60508 3388 60564 3390
rect 59052 1148 59108 1204
rect 70588 5964 70644 6020
rect 65660 5234 65716 5236
rect 65660 5182 65662 5234
rect 65662 5182 65714 5234
rect 65714 5182 65716 5234
rect 65660 5180 65716 5182
rect 63980 4844 64036 4900
rect 62188 2492 62244 2548
rect 62412 3442 62468 3444
rect 62412 3390 62414 3442
rect 62414 3390 62466 3442
rect 62466 3390 62468 3442
rect 62412 3388 62468 3390
rect 64316 4844 64372 4900
rect 64092 4508 64148 4564
rect 64428 3442 64484 3444
rect 64428 3390 64430 3442
rect 64430 3390 64482 3442
rect 64482 3390 64484 3442
rect 64428 3388 64484 3390
rect 64092 2604 64148 2660
rect 67228 924 67284 980
rect 67340 3388 67396 3444
rect 68908 3442 68964 3444
rect 68908 3390 68910 3442
rect 68910 3390 68962 3442
rect 68962 3390 68964 3442
rect 68908 3388 68964 3390
rect 68684 1372 68740 1428
rect 70700 4172 70756 4228
rect 82796 12236 82852 12292
rect 74852 11002 74908 11004
rect 74852 10950 74854 11002
rect 74854 10950 74906 11002
rect 74906 10950 74908 11002
rect 74852 10948 74908 10950
rect 74956 11002 75012 11004
rect 74956 10950 74958 11002
rect 74958 10950 75010 11002
rect 75010 10950 75012 11002
rect 74956 10948 75012 10950
rect 75060 11002 75116 11004
rect 75060 10950 75062 11002
rect 75062 10950 75114 11002
rect 75114 10950 75116 11002
rect 75060 10948 75116 10950
rect 74732 10444 74788 10500
rect 74508 5740 74564 5796
rect 73836 5068 73892 5124
rect 73388 4956 73444 5012
rect 72604 4396 72660 4452
rect 71820 4226 71876 4228
rect 71820 4174 71822 4226
rect 71822 4174 71874 4226
rect 71874 4174 71876 4226
rect 71820 4172 71876 4174
rect 72716 3836 72772 3892
rect 73500 4450 73556 4452
rect 73500 4398 73502 4450
rect 73502 4398 73554 4450
rect 73554 4398 73556 4450
rect 73500 4396 73556 4398
rect 73836 4396 73892 4452
rect 73388 3836 73444 3892
rect 79436 9548 79492 9604
rect 74852 9434 74908 9436
rect 74852 9382 74854 9434
rect 74854 9382 74906 9434
rect 74906 9382 74908 9434
rect 74852 9380 74908 9382
rect 74956 9434 75012 9436
rect 74956 9382 74958 9434
rect 74958 9382 75010 9434
rect 75010 9382 75012 9434
rect 74956 9380 75012 9382
rect 75060 9434 75116 9436
rect 75060 9382 75062 9434
rect 75062 9382 75114 9434
rect 75114 9382 75116 9434
rect 75060 9380 75116 9382
rect 75628 8764 75684 8820
rect 74852 7866 74908 7868
rect 74852 7814 74854 7866
rect 74854 7814 74906 7866
rect 74906 7814 74908 7866
rect 74852 7812 74908 7814
rect 74956 7866 75012 7868
rect 74956 7814 74958 7866
rect 74958 7814 75010 7866
rect 75010 7814 75012 7866
rect 74956 7812 75012 7814
rect 75060 7866 75116 7868
rect 75060 7814 75062 7866
rect 75062 7814 75114 7866
rect 75114 7814 75116 7866
rect 75060 7812 75116 7814
rect 74852 6298 74908 6300
rect 74852 6246 74854 6298
rect 74854 6246 74906 6298
rect 74906 6246 74908 6298
rect 74852 6244 74908 6246
rect 74956 6298 75012 6300
rect 74956 6246 74958 6298
rect 74958 6246 75010 6298
rect 75010 6246 75012 6298
rect 74956 6244 75012 6246
rect 75060 6298 75116 6300
rect 75060 6246 75062 6298
rect 75062 6246 75114 6298
rect 75114 6246 75116 6298
rect 75060 6244 75116 6246
rect 75404 5010 75460 5012
rect 75404 4958 75406 5010
rect 75406 4958 75458 5010
rect 75458 4958 75460 5010
rect 75404 4956 75460 4958
rect 74852 4730 74908 4732
rect 74852 4678 74854 4730
rect 74854 4678 74906 4730
rect 74906 4678 74908 4730
rect 74852 4676 74908 4678
rect 74956 4730 75012 4732
rect 74956 4678 74958 4730
rect 74958 4678 75010 4730
rect 75010 4678 75012 4730
rect 74956 4676 75012 4678
rect 75060 4730 75116 4732
rect 75060 4678 75062 4730
rect 75062 4678 75114 4730
rect 75114 4678 75116 4730
rect 75060 4676 75116 4678
rect 76188 7980 76244 8036
rect 75740 5794 75796 5796
rect 75740 5742 75742 5794
rect 75742 5742 75794 5794
rect 75794 5742 75796 5794
rect 75740 5740 75796 5742
rect 77980 7308 78036 7364
rect 76188 4956 76244 5012
rect 77196 5404 77252 5460
rect 75628 4450 75684 4452
rect 75628 4398 75630 4450
rect 75630 4398 75682 4450
rect 75682 4398 75684 4450
rect 75628 4396 75684 4398
rect 75740 3612 75796 3668
rect 73164 3330 73220 3332
rect 73164 3278 73166 3330
rect 73166 3278 73218 3330
rect 73218 3278 73220 3330
rect 73164 3276 73220 3278
rect 74852 3162 74908 3164
rect 74852 3110 74854 3162
rect 74854 3110 74906 3162
rect 74906 3110 74908 3162
rect 74852 3108 74908 3110
rect 74956 3162 75012 3164
rect 74956 3110 74958 3162
rect 74958 3110 75010 3162
rect 75010 3110 75012 3162
rect 74956 3108 75012 3110
rect 75060 3162 75116 3164
rect 75060 3110 75062 3162
rect 75062 3110 75114 3162
rect 75114 3110 75116 3162
rect 75060 3108 75116 3110
rect 77644 5404 77700 5460
rect 78540 5122 78596 5124
rect 78540 5070 78542 5122
rect 78542 5070 78594 5122
rect 78594 5070 78596 5122
rect 78540 5068 78596 5070
rect 76972 3666 77028 3668
rect 76972 3614 76974 3666
rect 76974 3614 77026 3666
rect 77026 3614 77028 3666
rect 76972 3612 77028 3614
rect 77420 3612 77476 3668
rect 78876 5068 78932 5124
rect 79436 5068 79492 5124
rect 79772 8988 79828 9044
rect 80668 8876 80724 8932
rect 80556 7420 80612 7476
rect 80556 5404 80612 5460
rect 98476 12124 98532 12180
rect 93262 11786 93318 11788
rect 93262 11734 93264 11786
rect 93264 11734 93316 11786
rect 93316 11734 93318 11786
rect 93262 11732 93318 11734
rect 93366 11786 93422 11788
rect 93366 11734 93368 11786
rect 93368 11734 93420 11786
rect 93420 11734 93422 11786
rect 93366 11732 93422 11734
rect 93470 11786 93526 11788
rect 93470 11734 93472 11786
rect 93472 11734 93524 11786
rect 93524 11734 93526 11786
rect 93470 11732 93526 11734
rect 98028 11116 98084 11172
rect 85596 10332 85652 10388
rect 81004 5122 81060 5124
rect 81004 5070 81006 5122
rect 81006 5070 81058 5122
rect 81058 5070 81060 5122
rect 81004 5068 81060 5070
rect 81452 5122 81508 5124
rect 81452 5070 81454 5122
rect 81454 5070 81506 5122
rect 81506 5070 81508 5122
rect 81452 5068 81508 5070
rect 82236 5122 82292 5124
rect 82236 5070 82238 5122
rect 82238 5070 82290 5122
rect 82290 5070 82292 5122
rect 82236 5068 82292 5070
rect 85372 6188 85428 6244
rect 82796 5068 82852 5124
rect 83356 5122 83412 5124
rect 83356 5070 83358 5122
rect 83358 5070 83410 5122
rect 83410 5070 83412 5122
rect 83356 5068 83412 5070
rect 83804 5122 83860 5124
rect 83804 5070 83806 5122
rect 83806 5070 83858 5122
rect 83858 5070 83860 5122
rect 83804 5068 83860 5070
rect 84588 5068 84644 5124
rect 78988 4172 79044 4228
rect 78988 3724 79044 3780
rect 78764 3666 78820 3668
rect 78764 3614 78766 3666
rect 78766 3614 78818 3666
rect 78818 3614 78820 3666
rect 78764 3612 78820 3614
rect 79100 3612 79156 3668
rect 80108 4338 80164 4340
rect 80108 4286 80110 4338
rect 80110 4286 80162 4338
rect 80162 4286 80164 4338
rect 80108 4284 80164 4286
rect 80556 4338 80612 4340
rect 80556 4286 80558 4338
rect 80558 4286 80610 4338
rect 80610 4286 80612 4338
rect 80556 4284 80612 4286
rect 81452 4338 81508 4340
rect 81452 4286 81454 4338
rect 81454 4286 81506 4338
rect 81506 4286 81508 4338
rect 81452 4284 81508 4286
rect 80780 3948 80836 4004
rect 80892 3666 80948 3668
rect 80892 3614 80894 3666
rect 80894 3614 80946 3666
rect 80946 3614 80948 3666
rect 80892 3612 80948 3614
rect 82124 4284 82180 4340
rect 83916 4844 83972 4900
rect 83020 4172 83076 4228
rect 82684 3948 82740 4004
rect 82124 2604 82180 2660
rect 82460 3388 82516 3444
rect 83356 3388 83412 3444
rect 85372 5068 85428 5124
rect 85484 5010 85540 5012
rect 85484 4958 85486 5010
rect 85486 4958 85538 5010
rect 85538 4958 85540 5010
rect 85484 4956 85540 4958
rect 83916 812 83972 868
rect 87164 10332 87220 10388
rect 86940 6130 86996 6132
rect 86940 6078 86942 6130
rect 86942 6078 86994 6130
rect 86994 6078 86996 6130
rect 86940 6076 86996 6078
rect 86044 5794 86100 5796
rect 86044 5742 86046 5794
rect 86046 5742 86098 5794
rect 86098 5742 86100 5794
rect 86044 5740 86100 5742
rect 86940 5740 86996 5796
rect 86044 4956 86100 5012
rect 86380 3948 86436 4004
rect 85596 3276 85652 3332
rect 85820 3836 85876 3892
rect 86716 3836 86772 3892
rect 93262 10218 93318 10220
rect 93262 10166 93264 10218
rect 93264 10166 93316 10218
rect 93316 10166 93318 10218
rect 93262 10164 93318 10166
rect 93366 10218 93422 10220
rect 93366 10166 93368 10218
rect 93368 10166 93420 10218
rect 93420 10166 93422 10218
rect 93366 10164 93422 10166
rect 93470 10218 93526 10220
rect 93470 10166 93472 10218
rect 93472 10166 93524 10218
rect 93524 10166 93526 10218
rect 93470 10164 93526 10166
rect 90748 9884 90804 9940
rect 90300 8876 90356 8932
rect 88396 6636 88452 6692
rect 87164 5180 87220 5236
rect 87836 6076 87892 6132
rect 87724 5010 87780 5012
rect 87724 4958 87726 5010
rect 87726 4958 87778 5010
rect 87778 4958 87780 5010
rect 87724 4956 87780 4958
rect 88396 6130 88452 6132
rect 88396 6078 88398 6130
rect 88398 6078 88450 6130
rect 88450 6078 88452 6130
rect 88396 6076 88452 6078
rect 88956 5852 89012 5908
rect 88172 4956 88228 5012
rect 89404 5180 89460 5236
rect 89852 5234 89908 5236
rect 89852 5182 89854 5234
rect 89854 5182 89906 5234
rect 89906 5182 89908 5234
rect 89852 5180 89908 5182
rect 90188 5180 90244 5236
rect 88956 4956 89012 5012
rect 87388 4060 87444 4116
rect 87500 3612 87556 3668
rect 86156 3330 86212 3332
rect 86156 3278 86158 3330
rect 86158 3278 86210 3330
rect 86210 3278 86212 3330
rect 86156 3276 86212 3278
rect 88284 4396 88340 4452
rect 89292 4450 89348 4452
rect 89292 4398 89294 4450
rect 89294 4398 89346 4450
rect 89346 4398 89348 4450
rect 89292 4396 89348 4398
rect 89068 3724 89124 3780
rect 88732 3666 88788 3668
rect 88732 3614 88734 3666
rect 88734 3614 88786 3666
rect 88786 3614 88788 3666
rect 88732 3612 88788 3614
rect 89180 3612 89236 3668
rect 93262 8650 93318 8652
rect 93262 8598 93264 8650
rect 93264 8598 93316 8650
rect 93316 8598 93318 8650
rect 93262 8596 93318 8598
rect 93366 8650 93422 8652
rect 93366 8598 93368 8650
rect 93368 8598 93420 8650
rect 93420 8598 93422 8650
rect 93366 8596 93422 8598
rect 93470 8650 93526 8652
rect 93470 8598 93472 8650
rect 93472 8598 93524 8650
rect 93524 8598 93526 8650
rect 93470 8596 93526 8598
rect 90748 5234 90804 5236
rect 90748 5182 90750 5234
rect 90750 5182 90802 5234
rect 90802 5182 90804 5234
rect 90748 5180 90804 5182
rect 91532 7196 91588 7252
rect 93262 7082 93318 7084
rect 93262 7030 93264 7082
rect 93264 7030 93316 7082
rect 93316 7030 93318 7082
rect 93262 7028 93318 7030
rect 93366 7082 93422 7084
rect 93366 7030 93368 7082
rect 93368 7030 93420 7082
rect 93420 7030 93422 7082
rect 93366 7028 93422 7030
rect 93470 7082 93526 7084
rect 93470 7030 93472 7082
rect 93472 7030 93524 7082
rect 93524 7030 93526 7082
rect 93470 7028 93526 7030
rect 97356 5964 97412 6020
rect 96460 5628 96516 5684
rect 93262 5514 93318 5516
rect 93262 5462 93264 5514
rect 93264 5462 93316 5514
rect 93316 5462 93318 5514
rect 93262 5460 93318 5462
rect 93366 5514 93422 5516
rect 93366 5462 93368 5514
rect 93368 5462 93420 5514
rect 93420 5462 93422 5514
rect 93366 5460 93422 5462
rect 93470 5514 93526 5516
rect 93470 5462 93472 5514
rect 93472 5462 93524 5514
rect 93524 5462 93526 5514
rect 93470 5460 93526 5462
rect 96460 5404 96516 5460
rect 96236 5346 96292 5348
rect 96236 5294 96238 5346
rect 96238 5294 96290 5346
rect 96290 5294 96292 5346
rect 96236 5292 96292 5294
rect 91532 4732 91588 4788
rect 94108 5180 94164 5236
rect 90300 4396 90356 4452
rect 90524 4450 90580 4452
rect 90524 4398 90526 4450
rect 90526 4398 90578 4450
rect 90578 4398 90580 4450
rect 90524 4396 90580 4398
rect 91084 4396 91140 4452
rect 93996 4450 94052 4452
rect 93996 4398 93998 4450
rect 93998 4398 94050 4450
rect 94050 4398 94052 4450
rect 93996 4396 94052 4398
rect 90860 4172 90916 4228
rect 90524 3666 90580 3668
rect 90524 3614 90526 3666
rect 90526 3614 90578 3666
rect 90578 3614 90580 3666
rect 90524 3612 90580 3614
rect 91756 4226 91812 4228
rect 91756 4174 91758 4226
rect 91758 4174 91810 4226
rect 91810 4174 91812 4226
rect 91756 4172 91812 4174
rect 93262 3946 93318 3948
rect 93262 3894 93264 3946
rect 93264 3894 93316 3946
rect 93316 3894 93318 3946
rect 93262 3892 93318 3894
rect 93366 3946 93422 3948
rect 93366 3894 93368 3946
rect 93368 3894 93420 3946
rect 93420 3894 93422 3946
rect 93366 3892 93422 3894
rect 93470 3946 93526 3948
rect 93470 3894 93472 3946
rect 93472 3894 93524 3946
rect 93524 3894 93526 3946
rect 93470 3892 93526 3894
rect 95452 5122 95508 5124
rect 95452 5070 95454 5122
rect 95454 5070 95506 5122
rect 95506 5070 95508 5122
rect 95452 5068 95508 5070
rect 94220 4396 94276 4452
rect 94556 4450 94612 4452
rect 94556 4398 94558 4450
rect 94558 4398 94610 4450
rect 94610 4398 94612 4450
rect 94556 4396 94612 4398
rect 97020 5404 97076 5460
rect 97916 6018 97972 6020
rect 97916 5966 97918 6018
rect 97918 5966 97970 6018
rect 97970 5966 97972 6018
rect 97916 5964 97972 5966
rect 97468 5628 97524 5684
rect 99036 5964 99092 6020
rect 97132 5068 97188 5124
rect 95228 3442 95284 3444
rect 95228 3390 95230 3442
rect 95230 3390 95282 3442
rect 95282 3390 95284 3442
rect 95228 3388 95284 3390
rect 95900 3388 95956 3444
rect 94668 1596 94724 1652
rect 96236 3442 96292 3444
rect 96236 3390 96238 3442
rect 96238 3390 96290 3442
rect 96290 3390 96292 3442
rect 96236 3388 96292 3390
rect 97580 3388 97636 3444
rect 99260 5122 99316 5124
rect 99260 5070 99262 5122
rect 99262 5070 99314 5122
rect 99314 5070 99316 5122
rect 99260 5068 99316 5070
rect 101164 12850 101220 12852
rect 101164 12798 101166 12850
rect 101166 12798 101218 12850
rect 101218 12798 101220 12850
rect 101164 12796 101220 12798
rect 101500 12850 101556 12852
rect 101500 12798 101502 12850
rect 101502 12798 101554 12850
rect 101554 12798 101556 12850
rect 101500 12796 101556 12798
rect 100156 12178 100212 12180
rect 100156 12126 100158 12178
rect 100158 12126 100210 12178
rect 100210 12126 100212 12178
rect 100156 12124 100212 12126
rect 100492 11170 100548 11172
rect 100492 11118 100494 11170
rect 100494 11118 100546 11170
rect 100546 11118 100548 11170
rect 100492 11116 100548 11118
rect 101164 11116 101220 11172
rect 101500 11170 101556 11172
rect 101500 11118 101502 11170
rect 101502 11118 101554 11170
rect 101554 11118 101556 11170
rect 101500 11116 101556 11118
rect 101948 10556 102004 10612
rect 101500 7644 101556 7700
rect 101948 5964 102004 6020
rect 102732 6018 102788 6020
rect 102732 5966 102734 6018
rect 102734 5966 102786 6018
rect 102786 5966 102788 6018
rect 102732 5964 102788 5966
rect 101164 5292 101220 5348
rect 101388 5852 101444 5908
rect 99484 5068 99540 5124
rect 98252 4172 98308 4228
rect 98588 4956 98644 5012
rect 98924 5010 98980 5012
rect 98924 4958 98926 5010
rect 98926 4958 98978 5010
rect 98978 4958 98980 5010
rect 98924 4956 98980 4958
rect 99036 4226 99092 4228
rect 99036 4174 99038 4226
rect 99038 4174 99090 4226
rect 99090 4174 99092 4226
rect 99036 4172 99092 4174
rect 101052 5122 101108 5124
rect 101052 5070 101054 5122
rect 101054 5070 101106 5122
rect 101106 5070 101108 5122
rect 101052 5068 101108 5070
rect 98028 3442 98084 3444
rect 98028 3390 98030 3442
rect 98030 3390 98082 3442
rect 98082 3390 98084 3442
rect 98028 3388 98084 3390
rect 99260 3388 99316 3444
rect 100828 3442 100884 3444
rect 100828 3390 100830 3442
rect 100830 3390 100882 3442
rect 100882 3390 100884 3442
rect 100828 3388 100884 3390
rect 102172 5852 102228 5908
rect 102620 5906 102676 5908
rect 102620 5854 102622 5906
rect 102622 5854 102674 5906
rect 102674 5854 102676 5906
rect 102620 5852 102676 5854
rect 105868 10780 105924 10836
rect 103740 5852 103796 5908
rect 101388 3724 101444 3780
rect 103292 3948 103348 4004
rect 103740 5292 103796 5348
rect 103852 5068 103908 5124
rect 103964 5010 104020 5012
rect 103964 4958 103966 5010
rect 103966 4958 104018 5010
rect 104018 4958 104020 5010
rect 103964 4956 104020 4958
rect 105532 7308 105588 7364
rect 106652 7308 106708 7364
rect 107772 15036 107828 15092
rect 105644 5180 105700 5236
rect 105868 5292 105924 5348
rect 104412 4956 104468 5012
rect 105644 4732 105700 4788
rect 104300 3948 104356 4004
rect 104300 3500 104356 3556
rect 101836 2268 101892 2324
rect 103068 3442 103124 3444
rect 103068 3390 103070 3442
rect 103070 3390 103122 3442
rect 103122 3390 103124 3442
rect 103068 3388 103124 3390
rect 104748 3442 104804 3444
rect 104748 3390 104750 3442
rect 104750 3390 104802 3442
rect 104802 3390 104804 3442
rect 104748 3388 104804 3390
rect 105980 3388 106036 3444
rect 106204 3500 106260 3556
rect 106316 3948 106372 4004
rect 109116 6748 109172 6804
rect 109116 6188 109172 6244
rect 109900 6188 109956 6244
rect 109788 5906 109844 5908
rect 109788 5854 109790 5906
rect 109790 5854 109842 5906
rect 109842 5854 109844 5906
rect 109788 5852 109844 5854
rect 107100 4732 107156 4788
rect 107436 3836 107492 3892
rect 106428 3612 106484 3668
rect 107660 3666 107716 3668
rect 107660 3614 107662 3666
rect 107662 3614 107714 3666
rect 107714 3614 107716 3666
rect 107660 3612 107716 3614
rect 106764 3554 106820 3556
rect 106764 3502 106766 3554
rect 106766 3502 106818 3554
rect 106818 3502 106820 3554
rect 106764 3500 106820 3502
rect 109564 5122 109620 5124
rect 109564 5070 109566 5122
rect 109566 5070 109618 5122
rect 109618 5070 109620 5122
rect 109564 5068 109620 5070
rect 111672 17274 111728 17276
rect 111672 17222 111674 17274
rect 111674 17222 111726 17274
rect 111726 17222 111728 17274
rect 111672 17220 111728 17222
rect 111776 17274 111832 17276
rect 111776 17222 111778 17274
rect 111778 17222 111830 17274
rect 111830 17222 111832 17274
rect 111776 17220 111832 17222
rect 111880 17274 111936 17276
rect 111880 17222 111882 17274
rect 111882 17222 111934 17274
rect 111934 17222 111936 17274
rect 111880 17220 111936 17222
rect 111672 15706 111728 15708
rect 111672 15654 111674 15706
rect 111674 15654 111726 15706
rect 111726 15654 111728 15706
rect 111672 15652 111728 15654
rect 111776 15706 111832 15708
rect 111776 15654 111778 15706
rect 111778 15654 111830 15706
rect 111830 15654 111832 15706
rect 111776 15652 111832 15654
rect 111880 15706 111936 15708
rect 111880 15654 111882 15706
rect 111882 15654 111934 15706
rect 111934 15654 111936 15706
rect 111880 15652 111936 15654
rect 111672 14138 111728 14140
rect 111672 14086 111674 14138
rect 111674 14086 111726 14138
rect 111726 14086 111728 14138
rect 111672 14084 111728 14086
rect 111776 14138 111832 14140
rect 111776 14086 111778 14138
rect 111778 14086 111830 14138
rect 111830 14086 111832 14138
rect 111776 14084 111832 14086
rect 111880 14138 111936 14140
rect 111880 14086 111882 14138
rect 111882 14086 111934 14138
rect 111934 14086 111936 14138
rect 111880 14084 111936 14086
rect 111672 12570 111728 12572
rect 111672 12518 111674 12570
rect 111674 12518 111726 12570
rect 111726 12518 111728 12570
rect 111672 12516 111728 12518
rect 111776 12570 111832 12572
rect 111776 12518 111778 12570
rect 111778 12518 111830 12570
rect 111830 12518 111832 12570
rect 111776 12516 111832 12518
rect 111880 12570 111936 12572
rect 111880 12518 111882 12570
rect 111882 12518 111934 12570
rect 111934 12518 111936 12570
rect 111880 12516 111936 12518
rect 111672 11002 111728 11004
rect 111672 10950 111674 11002
rect 111674 10950 111726 11002
rect 111726 10950 111728 11002
rect 111672 10948 111728 10950
rect 111776 11002 111832 11004
rect 111776 10950 111778 11002
rect 111778 10950 111830 11002
rect 111830 10950 111832 11002
rect 111776 10948 111832 10950
rect 111880 11002 111936 11004
rect 111880 10950 111882 11002
rect 111882 10950 111934 11002
rect 111934 10950 111936 11002
rect 111880 10948 111936 10950
rect 111672 9434 111728 9436
rect 111672 9382 111674 9434
rect 111674 9382 111726 9434
rect 111726 9382 111728 9434
rect 111672 9380 111728 9382
rect 111776 9434 111832 9436
rect 111776 9382 111778 9434
rect 111778 9382 111830 9434
rect 111830 9382 111832 9434
rect 111776 9380 111832 9382
rect 111880 9434 111936 9436
rect 111880 9382 111882 9434
rect 111882 9382 111934 9434
rect 111934 9382 111936 9434
rect 111880 9380 111936 9382
rect 111672 7866 111728 7868
rect 111672 7814 111674 7866
rect 111674 7814 111726 7866
rect 111726 7814 111728 7866
rect 111672 7812 111728 7814
rect 111776 7866 111832 7868
rect 111776 7814 111778 7866
rect 111778 7814 111830 7866
rect 111830 7814 111832 7866
rect 111776 7812 111832 7814
rect 111880 7866 111936 7868
rect 111880 7814 111882 7866
rect 111882 7814 111934 7866
rect 111934 7814 111936 7866
rect 111880 7812 111936 7814
rect 110460 5852 110516 5908
rect 109788 5068 109844 5124
rect 107884 3388 107940 3444
rect 108332 4844 108388 4900
rect 106092 2380 106148 2436
rect 109228 4508 109284 4564
rect 109564 3948 109620 4004
rect 109340 3612 109396 3668
rect 108668 3442 108724 3444
rect 108668 3390 108670 3442
rect 108670 3390 108722 3442
rect 108722 3390 108724 3442
rect 108668 3388 108724 3390
rect 108332 2492 108388 2548
rect 110908 4172 110964 4228
rect 111672 6298 111728 6300
rect 111672 6246 111674 6298
rect 111674 6246 111726 6298
rect 111726 6246 111728 6298
rect 111672 6244 111728 6246
rect 111776 6298 111832 6300
rect 111776 6246 111778 6298
rect 111778 6246 111830 6298
rect 111830 6246 111832 6298
rect 111776 6244 111832 6246
rect 111880 6298 111936 6300
rect 111880 6246 111882 6298
rect 111882 6246 111934 6298
rect 111934 6246 111936 6298
rect 111880 6244 111936 6246
rect 112028 5740 112084 5796
rect 111468 5122 111524 5124
rect 111468 5070 111470 5122
rect 111470 5070 111522 5122
rect 111522 5070 111524 5122
rect 111468 5068 111524 5070
rect 111020 3948 111076 4004
rect 110908 3612 110964 3668
rect 111020 3500 111076 3556
rect 110684 2492 110740 2548
rect 111672 4730 111728 4732
rect 111672 4678 111674 4730
rect 111674 4678 111726 4730
rect 111726 4678 111728 4730
rect 111672 4676 111728 4678
rect 111776 4730 111832 4732
rect 111776 4678 111778 4730
rect 111778 4678 111830 4730
rect 111830 4678 111832 4730
rect 111776 4676 111832 4678
rect 111880 4730 111936 4732
rect 111880 4678 111882 4730
rect 111882 4678 111934 4730
rect 111934 4678 111936 4730
rect 111880 4676 111936 4678
rect 111804 4226 111860 4228
rect 111804 4174 111806 4226
rect 111806 4174 111858 4226
rect 111858 4174 111860 4226
rect 111804 4172 111860 4174
rect 114268 20524 114324 20580
rect 114268 18620 114324 18676
rect 115836 18284 115892 18340
rect 115836 15036 115892 15092
rect 117404 14364 117460 14420
rect 115276 9100 115332 9156
rect 115276 5964 115332 6020
rect 116060 6018 116116 6020
rect 116060 5966 116062 6018
rect 116062 5966 116114 6018
rect 116114 5966 116116 6018
rect 116060 5964 116116 5966
rect 115388 5852 115444 5908
rect 113148 5122 113204 5124
rect 113148 5070 113150 5122
rect 113150 5070 113202 5122
rect 113202 5070 113204 5122
rect 113148 5068 113204 5070
rect 111672 3162 111728 3164
rect 111672 3110 111674 3162
rect 111674 3110 111726 3162
rect 111726 3110 111728 3162
rect 111672 3108 111728 3110
rect 111776 3162 111832 3164
rect 111776 3110 111778 3162
rect 111778 3110 111830 3162
rect 111830 3110 111832 3162
rect 111776 3108 111832 3110
rect 111880 3162 111936 3164
rect 111880 3110 111882 3162
rect 111882 3110 111934 3162
rect 111934 3110 111936 3162
rect 111880 3108 111936 3110
rect 111132 2828 111188 2884
rect 112588 3500 112644 3556
rect 112700 3388 112756 3444
rect 112252 2828 112308 2884
rect 117964 7532 118020 7588
rect 119196 6748 119252 6804
rect 119308 6972 119364 7028
rect 116508 6018 116564 6020
rect 116508 5966 116510 6018
rect 116510 5966 116562 6018
rect 116562 5966 116564 6018
rect 116508 5964 116564 5966
rect 117740 5964 117796 6020
rect 113820 4172 113876 4228
rect 114380 4226 114436 4228
rect 114380 4174 114382 4226
rect 114382 4174 114434 4226
rect 114434 4174 114436 4226
rect 114380 4172 114436 4174
rect 113484 3554 113540 3556
rect 113484 3502 113486 3554
rect 113486 3502 113538 3554
rect 113538 3502 113540 3554
rect 113484 3500 113540 3502
rect 113260 3388 113316 3444
rect 113932 3442 113988 3444
rect 113932 3390 113934 3442
rect 113934 3390 113986 3442
rect 113986 3390 113988 3442
rect 113932 3388 113988 3390
rect 114828 3442 114884 3444
rect 114828 3390 114830 3442
rect 114830 3390 114882 3442
rect 114882 3390 114884 3442
rect 114828 3388 114884 3390
rect 113036 1036 113092 1092
rect 115724 4956 115780 5012
rect 115388 4226 115444 4228
rect 115388 4174 115390 4226
rect 115390 4174 115442 4226
rect 115442 4174 115444 4226
rect 115388 4172 115444 4174
rect 115612 3442 115668 3444
rect 115612 3390 115614 3442
rect 115614 3390 115666 3442
rect 115666 3390 115668 3442
rect 115612 3388 115668 3390
rect 115836 3612 115892 3668
rect 116060 4172 116116 4228
rect 115724 2716 115780 2772
rect 115052 1484 115108 1540
rect 117180 5010 117236 5012
rect 117180 4958 117182 5010
rect 117182 4958 117234 5010
rect 117234 4958 117236 5010
rect 117180 4956 117236 4958
rect 119084 5906 119140 5908
rect 119084 5854 119086 5906
rect 119086 5854 119138 5906
rect 119138 5854 119140 5906
rect 119084 5852 119140 5854
rect 117068 4844 117124 4900
rect 116732 4172 116788 4228
rect 117516 4226 117572 4228
rect 117516 4174 117518 4226
rect 117518 4174 117570 4226
rect 117570 4174 117572 4226
rect 117516 4172 117572 4174
rect 116732 3666 116788 3668
rect 116732 3614 116734 3666
rect 116734 3614 116786 3666
rect 116786 3614 116788 3666
rect 116732 3612 116788 3614
rect 118300 5010 118356 5012
rect 118300 4958 118302 5010
rect 118302 4958 118354 5010
rect 118354 4958 118356 5010
rect 118300 4956 118356 4958
rect 118076 3836 118132 3892
rect 121772 23660 121828 23716
rect 121772 6972 121828 7028
rect 122108 10668 122164 10724
rect 120204 6748 120260 6804
rect 119756 5906 119812 5908
rect 119756 5854 119758 5906
rect 119758 5854 119810 5906
rect 119810 5854 119812 5906
rect 119756 5852 119812 5854
rect 119868 5010 119924 5012
rect 119868 4958 119870 5010
rect 119870 4958 119922 5010
rect 119922 4958 119924 5010
rect 119868 4956 119924 4958
rect 122668 7756 122724 7812
rect 122668 6076 122724 6132
rect 122108 5964 122164 6020
rect 122892 6018 122948 6020
rect 122892 5966 122894 6018
rect 122894 5966 122946 6018
rect 122946 5966 122948 6018
rect 122892 5964 122948 5966
rect 123900 5906 123956 5908
rect 123900 5854 123902 5906
rect 123902 5854 123954 5906
rect 123954 5854 123956 5906
rect 123900 5852 123956 5854
rect 123340 5740 123396 5796
rect 122332 5180 122388 5236
rect 123452 5180 123508 5236
rect 118972 4844 119028 4900
rect 120204 4562 120260 4564
rect 120204 4510 120206 4562
rect 120206 4510 120258 4562
rect 120258 4510 120260 4562
rect 120204 4508 120260 4510
rect 118748 3612 118804 3668
rect 117740 3388 117796 3444
rect 118524 3442 118580 3444
rect 118524 3390 118526 3442
rect 118526 3390 118578 3442
rect 118578 3390 118580 3442
rect 118524 3388 118580 3390
rect 120204 3836 120260 3892
rect 119644 3666 119700 3668
rect 119644 3614 119646 3666
rect 119646 3614 119698 3666
rect 119698 3614 119700 3666
rect 119644 3612 119700 3614
rect 120652 3612 120708 3668
rect 119196 3388 119252 3444
rect 119420 3388 119476 3444
rect 120652 3442 120708 3444
rect 120652 3390 120654 3442
rect 120654 3390 120706 3442
rect 120706 3390 120708 3442
rect 120652 3388 120708 3390
rect 121100 3388 121156 3444
rect 123116 5010 123172 5012
rect 123116 4958 123118 5010
rect 123118 4958 123170 5010
rect 123170 4958 123172 5010
rect 123116 4956 123172 4958
rect 121548 3666 121604 3668
rect 121548 3614 121550 3666
rect 121550 3614 121602 3666
rect 121602 3614 121604 3666
rect 121548 3612 121604 3614
rect 123788 5010 123844 5012
rect 123788 4958 123790 5010
rect 123790 4958 123842 5010
rect 123842 4958 123844 5010
rect 123788 4956 123844 4958
rect 126028 22876 126084 22932
rect 126924 8428 126980 8484
rect 124572 5906 124628 5908
rect 124572 5854 124574 5906
rect 124574 5854 124626 5906
rect 124626 5854 124628 5906
rect 124572 5852 124628 5854
rect 124348 5740 124404 5796
rect 125468 5740 125524 5796
rect 126588 5794 126644 5796
rect 126588 5742 126590 5794
rect 126590 5742 126642 5794
rect 126642 5742 126644 5794
rect 126588 5740 126644 5742
rect 124908 4956 124964 5012
rect 121436 3388 121492 3444
rect 121996 3442 122052 3444
rect 121996 3390 121998 3442
rect 121998 3390 122050 3442
rect 122050 3390 122052 3442
rect 121996 3388 122052 3390
rect 122780 3388 122836 3444
rect 121324 1260 121380 1316
rect 124348 3442 124404 3444
rect 124348 3390 124350 3442
rect 124350 3390 124402 3442
rect 124402 3390 124404 3442
rect 124348 3388 124404 3390
rect 125132 5010 125188 5012
rect 125132 4958 125134 5010
rect 125134 4958 125186 5010
rect 125186 4958 125188 5010
rect 125132 4956 125188 4958
rect 126812 5010 126868 5012
rect 126812 4958 126814 5010
rect 126814 4958 126866 5010
rect 126866 4958 126868 5010
rect 126812 4956 126868 4958
rect 127596 4620 127652 4676
rect 126812 4338 126868 4340
rect 126812 4286 126814 4338
rect 126814 4286 126866 4338
rect 126866 4286 126868 4338
rect 126812 4284 126868 4286
rect 130082 29034 130138 29036
rect 130082 28982 130084 29034
rect 130084 28982 130136 29034
rect 130136 28982 130138 29034
rect 130082 28980 130138 28982
rect 130186 29034 130242 29036
rect 130186 28982 130188 29034
rect 130188 28982 130240 29034
rect 130240 28982 130242 29034
rect 130186 28980 130242 28982
rect 130290 29034 130346 29036
rect 130290 28982 130292 29034
rect 130292 28982 130344 29034
rect 130344 28982 130346 29034
rect 130290 28980 130346 28982
rect 130082 27466 130138 27468
rect 130082 27414 130084 27466
rect 130084 27414 130136 27466
rect 130136 27414 130138 27466
rect 130082 27412 130138 27414
rect 130186 27466 130242 27468
rect 130186 27414 130188 27466
rect 130188 27414 130240 27466
rect 130240 27414 130242 27466
rect 130186 27412 130242 27414
rect 130290 27466 130346 27468
rect 130290 27414 130292 27466
rect 130292 27414 130344 27466
rect 130344 27414 130346 27466
rect 130290 27412 130346 27414
rect 130082 25898 130138 25900
rect 130082 25846 130084 25898
rect 130084 25846 130136 25898
rect 130136 25846 130138 25898
rect 130082 25844 130138 25846
rect 130186 25898 130242 25900
rect 130186 25846 130188 25898
rect 130188 25846 130240 25898
rect 130240 25846 130242 25898
rect 130186 25844 130242 25846
rect 130290 25898 130346 25900
rect 130290 25846 130292 25898
rect 130292 25846 130344 25898
rect 130344 25846 130346 25898
rect 130290 25844 130346 25846
rect 130082 24330 130138 24332
rect 130082 24278 130084 24330
rect 130084 24278 130136 24330
rect 130136 24278 130138 24330
rect 130082 24276 130138 24278
rect 130186 24330 130242 24332
rect 130186 24278 130188 24330
rect 130188 24278 130240 24330
rect 130240 24278 130242 24330
rect 130186 24276 130242 24278
rect 130290 24330 130346 24332
rect 130290 24278 130292 24330
rect 130292 24278 130344 24330
rect 130344 24278 130346 24330
rect 130290 24276 130346 24278
rect 130082 22762 130138 22764
rect 130082 22710 130084 22762
rect 130084 22710 130136 22762
rect 130136 22710 130138 22762
rect 130082 22708 130138 22710
rect 130186 22762 130242 22764
rect 130186 22710 130188 22762
rect 130188 22710 130240 22762
rect 130240 22710 130242 22762
rect 130186 22708 130242 22710
rect 130290 22762 130346 22764
rect 130290 22710 130292 22762
rect 130292 22710 130344 22762
rect 130344 22710 130346 22762
rect 130290 22708 130346 22710
rect 130082 21194 130138 21196
rect 130082 21142 130084 21194
rect 130084 21142 130136 21194
rect 130136 21142 130138 21194
rect 130082 21140 130138 21142
rect 130186 21194 130242 21196
rect 130186 21142 130188 21194
rect 130188 21142 130240 21194
rect 130240 21142 130242 21194
rect 130186 21140 130242 21142
rect 130290 21194 130346 21196
rect 130290 21142 130292 21194
rect 130292 21142 130344 21194
rect 130344 21142 130346 21194
rect 130290 21140 130346 21142
rect 130082 19626 130138 19628
rect 130082 19574 130084 19626
rect 130084 19574 130136 19626
rect 130136 19574 130138 19626
rect 130082 19572 130138 19574
rect 130186 19626 130242 19628
rect 130186 19574 130188 19626
rect 130188 19574 130240 19626
rect 130240 19574 130242 19626
rect 130186 19572 130242 19574
rect 130290 19626 130346 19628
rect 130290 19574 130292 19626
rect 130292 19574 130344 19626
rect 130344 19574 130346 19626
rect 130290 19572 130346 19574
rect 130082 18058 130138 18060
rect 130082 18006 130084 18058
rect 130084 18006 130136 18058
rect 130136 18006 130138 18058
rect 130082 18004 130138 18006
rect 130186 18058 130242 18060
rect 130186 18006 130188 18058
rect 130188 18006 130240 18058
rect 130240 18006 130242 18058
rect 130186 18004 130242 18006
rect 130290 18058 130346 18060
rect 130290 18006 130292 18058
rect 130292 18006 130344 18058
rect 130344 18006 130346 18058
rect 130290 18004 130346 18006
rect 130082 16490 130138 16492
rect 130082 16438 130084 16490
rect 130084 16438 130136 16490
rect 130136 16438 130138 16490
rect 130082 16436 130138 16438
rect 130186 16490 130242 16492
rect 130186 16438 130188 16490
rect 130188 16438 130240 16490
rect 130240 16438 130242 16490
rect 130186 16436 130242 16438
rect 130290 16490 130346 16492
rect 130290 16438 130292 16490
rect 130292 16438 130344 16490
rect 130344 16438 130346 16490
rect 130290 16436 130346 16438
rect 130082 14922 130138 14924
rect 130082 14870 130084 14922
rect 130084 14870 130136 14922
rect 130136 14870 130138 14922
rect 130082 14868 130138 14870
rect 130186 14922 130242 14924
rect 130186 14870 130188 14922
rect 130188 14870 130240 14922
rect 130240 14870 130242 14922
rect 130186 14868 130242 14870
rect 130290 14922 130346 14924
rect 130290 14870 130292 14922
rect 130292 14870 130344 14922
rect 130344 14870 130346 14922
rect 130290 14868 130346 14870
rect 130508 14140 130564 14196
rect 130082 13354 130138 13356
rect 130082 13302 130084 13354
rect 130084 13302 130136 13354
rect 130136 13302 130138 13354
rect 130082 13300 130138 13302
rect 130186 13354 130242 13356
rect 130186 13302 130188 13354
rect 130188 13302 130240 13354
rect 130240 13302 130242 13354
rect 130186 13300 130242 13302
rect 130290 13354 130346 13356
rect 130290 13302 130292 13354
rect 130292 13302 130344 13354
rect 130344 13302 130346 13354
rect 130290 13300 130346 13302
rect 130082 11786 130138 11788
rect 130082 11734 130084 11786
rect 130084 11734 130136 11786
rect 130136 11734 130138 11786
rect 130082 11732 130138 11734
rect 130186 11786 130242 11788
rect 130186 11734 130188 11786
rect 130188 11734 130240 11786
rect 130240 11734 130242 11786
rect 130186 11732 130242 11734
rect 130290 11786 130346 11788
rect 130290 11734 130292 11786
rect 130292 11734 130344 11786
rect 130344 11734 130346 11786
rect 130290 11732 130346 11734
rect 130082 10218 130138 10220
rect 130082 10166 130084 10218
rect 130084 10166 130136 10218
rect 130136 10166 130138 10218
rect 130082 10164 130138 10166
rect 130186 10218 130242 10220
rect 130186 10166 130188 10218
rect 130188 10166 130240 10218
rect 130240 10166 130242 10218
rect 130186 10164 130242 10166
rect 130290 10218 130346 10220
rect 130290 10166 130292 10218
rect 130292 10166 130344 10218
rect 130344 10166 130346 10218
rect 130290 10164 130346 10166
rect 130082 8650 130138 8652
rect 130082 8598 130084 8650
rect 130084 8598 130136 8650
rect 130136 8598 130138 8650
rect 130082 8596 130138 8598
rect 130186 8650 130242 8652
rect 130186 8598 130188 8650
rect 130188 8598 130240 8650
rect 130240 8598 130242 8650
rect 130186 8596 130242 8598
rect 130290 8650 130346 8652
rect 130290 8598 130292 8650
rect 130292 8598 130344 8650
rect 130344 8598 130346 8650
rect 130290 8596 130346 8598
rect 129836 7586 129892 7588
rect 129836 7534 129838 7586
rect 129838 7534 129890 7586
rect 129890 7534 129892 7586
rect 129836 7532 129892 7534
rect 128828 6860 128884 6916
rect 130082 7082 130138 7084
rect 130082 7030 130084 7082
rect 130084 7030 130136 7082
rect 130136 7030 130138 7082
rect 130082 7028 130138 7030
rect 130186 7082 130242 7084
rect 130186 7030 130188 7082
rect 130188 7030 130240 7082
rect 130240 7030 130242 7082
rect 130186 7028 130242 7030
rect 130290 7082 130346 7084
rect 130290 7030 130292 7082
rect 130292 7030 130344 7082
rect 130344 7030 130346 7082
rect 130290 7028 130346 7030
rect 128828 5964 128884 6020
rect 128940 5740 128996 5796
rect 127932 4620 127988 4676
rect 127820 4396 127876 4452
rect 127596 4114 127652 4116
rect 127596 4062 127598 4114
rect 127598 4062 127650 4114
rect 127650 4062 127652 4114
rect 127596 4060 127652 4062
rect 126140 3388 126196 3444
rect 124908 2940 124964 2996
rect 127372 3442 127428 3444
rect 127372 3390 127374 3442
rect 127374 3390 127426 3442
rect 127426 3390 127428 3442
rect 127372 3388 127428 3390
rect 128492 4060 128548 4116
rect 129500 6018 129556 6020
rect 129500 5966 129502 6018
rect 129502 5966 129554 6018
rect 129554 5966 129556 6018
rect 129500 5964 129556 5966
rect 130508 6130 130564 6132
rect 130508 6078 130510 6130
rect 130510 6078 130562 6130
rect 130562 6078 130564 6130
rect 130508 6076 130564 6078
rect 129948 5740 130004 5796
rect 130082 5514 130138 5516
rect 130082 5462 130084 5514
rect 130084 5462 130136 5514
rect 130136 5462 130138 5514
rect 130082 5460 130138 5462
rect 130186 5514 130242 5516
rect 130186 5462 130188 5514
rect 130188 5462 130240 5514
rect 130240 5462 130242 5514
rect 130186 5460 130242 5462
rect 130290 5514 130346 5516
rect 130290 5462 130292 5514
rect 130292 5462 130344 5514
rect 130344 5462 130346 5514
rect 130290 5460 130346 5462
rect 129276 4508 129332 4564
rect 129164 4450 129220 4452
rect 129164 4398 129166 4450
rect 129166 4398 129218 4450
rect 129218 4398 129220 4450
rect 129164 4396 129220 4398
rect 129276 4284 129332 4340
rect 130082 3946 130138 3948
rect 130082 3894 130084 3946
rect 130084 3894 130136 3946
rect 130136 3894 130138 3946
rect 130082 3892 130138 3894
rect 130186 3946 130242 3948
rect 130186 3894 130188 3946
rect 130188 3894 130240 3946
rect 130240 3894 130242 3946
rect 130186 3892 130242 3894
rect 130290 3946 130346 3948
rect 130290 3894 130292 3946
rect 130292 3894 130344 3946
rect 130344 3894 130346 3946
rect 130290 3892 130346 3894
rect 129276 3666 129332 3668
rect 129276 3614 129278 3666
rect 129278 3614 129330 3666
rect 129330 3614 129332 3666
rect 129276 3612 129332 3614
rect 129836 3666 129892 3668
rect 129836 3614 129838 3666
rect 129838 3614 129890 3666
rect 129890 3614 129892 3666
rect 129836 3612 129892 3614
rect 130620 4732 130676 4788
rect 131292 7586 131348 7588
rect 131292 7534 131294 7586
rect 131294 7534 131346 7586
rect 131346 7534 131348 7586
rect 131292 7532 131348 7534
rect 131964 11900 132020 11956
rect 131740 7586 131796 7588
rect 131740 7534 131742 7586
rect 131742 7534 131794 7586
rect 131794 7534 131796 7586
rect 131740 7532 131796 7534
rect 131068 6076 131124 6132
rect 130956 5740 131012 5796
rect 132636 5906 132692 5908
rect 132636 5854 132638 5906
rect 132638 5854 132690 5906
rect 132690 5854 132692 5906
rect 132636 5852 132692 5854
rect 132076 5740 132132 5796
rect 131740 5346 131796 5348
rect 131740 5294 131742 5346
rect 131742 5294 131794 5346
rect 131794 5294 131796 5346
rect 131740 5292 131796 5294
rect 130844 4956 130900 5012
rect 130508 3612 130564 3668
rect 128828 1148 128884 1204
rect 129500 3500 129556 3556
rect 133532 12012 133588 12068
rect 133532 7644 133588 7700
rect 133980 10332 134036 10388
rect 133644 6412 133700 6468
rect 132972 5292 133028 5348
rect 132972 5010 133028 5012
rect 132972 4958 132974 5010
rect 132974 4958 133026 5010
rect 133026 4958 133028 5010
rect 132972 4956 133028 4958
rect 133532 5122 133588 5124
rect 133532 5070 133534 5122
rect 133534 5070 133586 5122
rect 133586 5070 133588 5122
rect 133532 5068 133588 5070
rect 133308 4956 133364 5012
rect 132300 4172 132356 4228
rect 131180 3666 131236 3668
rect 131180 3614 131182 3666
rect 131182 3614 131234 3666
rect 131234 3614 131236 3666
rect 131180 3612 131236 3614
rect 132188 3500 132244 3556
rect 131180 3388 131236 3444
rect 132412 3388 132468 3444
rect 132860 4396 132916 4452
rect 133420 4226 133476 4228
rect 133420 4174 133422 4226
rect 133422 4174 133474 4226
rect 133474 4174 133476 4226
rect 133420 4172 133476 4174
rect 133756 5794 133812 5796
rect 133756 5742 133758 5794
rect 133758 5742 133810 5794
rect 133810 5742 133812 5794
rect 133756 5740 133812 5742
rect 136220 8764 136276 8820
rect 137004 6466 137060 6468
rect 137004 6414 137006 6466
rect 137006 6414 137058 6466
rect 137058 6414 137060 6466
rect 137004 6412 137060 6414
rect 136220 6130 136276 6132
rect 136220 6078 136222 6130
rect 136222 6078 136274 6130
rect 136274 6078 136276 6130
rect 136220 6076 136276 6078
rect 138572 29932 138628 29988
rect 138572 14140 138628 14196
rect 137564 10444 137620 10500
rect 142156 36258 142212 36260
rect 142156 36206 142158 36258
rect 142158 36206 142210 36258
rect 142210 36206 142212 36258
rect 142156 36204 142212 36206
rect 143052 36204 143108 36260
rect 144172 36316 144228 36372
rect 142156 35532 142212 35588
rect 141260 34636 141316 34692
rect 141036 28588 141092 28644
rect 139468 22988 139524 23044
rect 141036 22876 141092 22932
rect 139468 14364 139524 14420
rect 140028 12348 140084 12404
rect 139916 7698 139972 7700
rect 139916 7646 139918 7698
rect 139918 7646 139970 7698
rect 139970 7646 139972 7698
rect 139916 7644 139972 7646
rect 137564 6524 137620 6580
rect 138124 6578 138180 6580
rect 138124 6526 138126 6578
rect 138126 6526 138178 6578
rect 138178 6526 138180 6578
rect 138124 6524 138180 6526
rect 137788 6412 137844 6468
rect 138908 6524 138964 6580
rect 138684 6412 138740 6468
rect 138236 6076 138292 6132
rect 139692 6076 139748 6132
rect 138684 6018 138740 6020
rect 138684 5966 138686 6018
rect 138686 5966 138738 6018
rect 138738 5966 138740 6018
rect 138684 5964 138740 5966
rect 140364 5964 140420 6020
rect 134428 5906 134484 5908
rect 134428 5854 134430 5906
rect 134430 5854 134482 5906
rect 134482 5854 134484 5906
rect 134428 5852 134484 5854
rect 135436 5346 135492 5348
rect 135436 5294 135438 5346
rect 135438 5294 135490 5346
rect 135490 5294 135492 5346
rect 135436 5292 135492 5294
rect 134652 5122 134708 5124
rect 134652 5070 134654 5122
rect 134654 5070 134706 5122
rect 134706 5070 134708 5122
rect 134652 5068 134708 5070
rect 134428 4450 134484 4452
rect 134428 4398 134430 4450
rect 134430 4398 134482 4450
rect 134482 4398 134484 4450
rect 134428 4396 134484 4398
rect 133644 3836 133700 3892
rect 138908 5682 138964 5684
rect 138908 5630 138910 5682
rect 138910 5630 138962 5682
rect 138962 5630 138964 5682
rect 138908 5628 138964 5630
rect 137004 5292 137060 5348
rect 137340 5404 137396 5460
rect 139244 5346 139300 5348
rect 139244 5294 139246 5346
rect 139246 5294 139298 5346
rect 139298 5294 139300 5346
rect 139244 5292 139300 5294
rect 136556 5122 136612 5124
rect 136556 5070 136558 5122
rect 136558 5070 136610 5122
rect 136610 5070 136612 5122
rect 136556 5068 136612 5070
rect 135884 4956 135940 5012
rect 136444 5010 136500 5012
rect 136444 4958 136446 5010
rect 136446 4958 136498 5010
rect 136498 4958 136500 5010
rect 136444 4956 136500 4958
rect 135772 4450 135828 4452
rect 135772 4398 135774 4450
rect 135774 4398 135826 4450
rect 135826 4398 135828 4450
rect 135772 4396 135828 4398
rect 135324 3500 135380 3556
rect 134204 3442 134260 3444
rect 134204 3390 134206 3442
rect 134206 3390 134258 3442
rect 134258 3390 134260 3442
rect 134204 3388 134260 3390
rect 134540 3388 134596 3444
rect 136108 3442 136164 3444
rect 136108 3390 136110 3442
rect 136110 3390 136162 3442
rect 136162 3390 136164 3442
rect 136108 3388 136164 3390
rect 136220 3500 136276 3556
rect 137004 3554 137060 3556
rect 137004 3502 137006 3554
rect 137006 3502 137058 3554
rect 137058 3502 137060 3554
rect 137004 3500 137060 3502
rect 138460 5122 138516 5124
rect 138460 5070 138462 5122
rect 138462 5070 138514 5122
rect 138514 5070 138516 5122
rect 138460 5068 138516 5070
rect 138348 5010 138404 5012
rect 138348 4958 138350 5010
rect 138350 4958 138402 5010
rect 138402 4958 138404 5010
rect 138348 4956 138404 4958
rect 138012 3388 138068 3444
rect 138124 4172 138180 4228
rect 138236 3330 138292 3332
rect 138236 3278 138238 3330
rect 138238 3278 138290 3330
rect 138290 3278 138292 3330
rect 138236 3276 138292 3278
rect 136444 924 136500 980
rect 139804 4956 139860 5012
rect 139020 4226 139076 4228
rect 139020 4174 139022 4226
rect 139022 4174 139074 4226
rect 139074 4174 139076 4226
rect 139020 4172 139076 4174
rect 140028 4172 140084 4228
rect 138348 1372 138404 1428
rect 139580 3388 139636 3444
rect 141148 6130 141204 6132
rect 141148 6078 141150 6130
rect 141150 6078 141202 6130
rect 141202 6078 141204 6130
rect 141148 6076 141204 6078
rect 144844 36316 144900 36372
rect 145964 36204 146020 36260
rect 143500 21420 143556 21476
rect 142716 9548 142772 9604
rect 142716 7980 142772 8036
rect 140924 5404 140980 5460
rect 143164 6524 143220 6580
rect 141820 5292 141876 5348
rect 142940 5628 142996 5684
rect 141148 5122 141204 5124
rect 141148 5070 141150 5122
rect 141150 5070 141202 5122
rect 141202 5070 141204 5122
rect 141148 5068 141204 5070
rect 140812 4172 140868 4228
rect 142156 4396 142212 4452
rect 141820 4226 141876 4228
rect 141820 4174 141822 4226
rect 141822 4174 141874 4226
rect 141874 4174 141876 4226
rect 141820 4172 141876 4174
rect 142044 4172 142100 4228
rect 141148 3724 141204 3780
rect 141484 3724 141540 3780
rect 140140 3388 140196 3444
rect 140924 3442 140980 3444
rect 140924 3390 140926 3442
rect 140926 3390 140978 3442
rect 140978 3390 140980 3442
rect 140924 3388 140980 3390
rect 141260 3388 141316 3444
rect 141820 3442 141876 3444
rect 141820 3390 141822 3442
rect 141822 3390 141874 3442
rect 141874 3390 141876 3442
rect 141820 3388 141876 3390
rect 143500 5852 143556 5908
rect 143948 18956 144004 19012
rect 143836 4450 143892 4452
rect 143836 4398 143838 4450
rect 143838 4398 143890 4450
rect 143890 4398 143892 4450
rect 143836 4396 143892 4398
rect 142716 3388 142772 3444
rect 142940 3388 142996 3444
rect 142044 2604 142100 2660
rect 144060 5740 144116 5796
rect 144284 35586 144340 35588
rect 144284 35534 144286 35586
rect 144286 35534 144338 35586
rect 144338 35534 144340 35586
rect 144284 35532 144340 35534
rect 144956 35532 145012 35588
rect 146076 35196 146132 35252
rect 144396 34690 144452 34692
rect 144396 34638 144398 34690
rect 144398 34638 144450 34690
rect 144450 34638 144452 34690
rect 144396 34636 144452 34638
rect 144956 34636 145012 34692
rect 146636 34690 146692 34692
rect 146636 34638 146638 34690
rect 146638 34638 146690 34690
rect 146690 34638 146692 34690
rect 146636 34636 146692 34638
rect 147756 36988 147812 37044
rect 148492 36090 148548 36092
rect 148492 36038 148494 36090
rect 148494 36038 148546 36090
rect 148546 36038 148548 36090
rect 148492 36036 148548 36038
rect 148596 36090 148652 36092
rect 148596 36038 148598 36090
rect 148598 36038 148650 36090
rect 148650 36038 148652 36090
rect 148596 36036 148652 36038
rect 148700 36090 148756 36092
rect 148700 36038 148702 36090
rect 148702 36038 148754 36090
rect 148754 36038 148756 36090
rect 148700 36036 148756 36038
rect 146076 34300 146132 34356
rect 144284 34018 144340 34020
rect 144284 33966 144286 34018
rect 144286 33966 144338 34018
rect 144338 33966 144340 34018
rect 144284 33964 144340 33966
rect 144956 33964 145012 34020
rect 146076 33404 146132 33460
rect 144396 33122 144452 33124
rect 144396 33070 144398 33122
rect 144398 33070 144450 33122
rect 144450 33070 144452 33122
rect 144396 33068 144452 33070
rect 144956 33068 145012 33124
rect 146076 32508 146132 32564
rect 144396 31554 144452 31556
rect 144396 31502 144398 31554
rect 144398 31502 144450 31554
rect 144450 31502 144452 31554
rect 144396 31500 144452 31502
rect 146076 31666 146132 31668
rect 146076 31614 146078 31666
rect 146078 31614 146130 31666
rect 146130 31614 146132 31666
rect 146076 31612 146132 31614
rect 144956 31500 145012 31556
rect 144284 30882 144340 30884
rect 144284 30830 144286 30882
rect 144286 30830 144338 30882
rect 144338 30830 144340 30882
rect 144284 30828 144340 30830
rect 144956 30828 145012 30884
rect 146076 30716 146132 30772
rect 144396 29986 144452 29988
rect 144396 29934 144398 29986
rect 144398 29934 144450 29986
rect 144450 29934 144452 29986
rect 144396 29932 144452 29934
rect 144956 29932 145012 29988
rect 146076 29932 146132 29988
rect 144284 29314 144340 29316
rect 144284 29262 144286 29314
rect 144286 29262 144338 29314
rect 144338 29262 144340 29314
rect 144284 29260 144340 29262
rect 144956 29260 145012 29316
rect 146076 28924 146132 28980
rect 144396 28642 144452 28644
rect 144396 28590 144398 28642
rect 144398 28590 144450 28642
rect 144450 28590 144452 28642
rect 144396 28588 144452 28590
rect 144956 28642 145012 28644
rect 144956 28590 144958 28642
rect 144958 28590 145010 28642
rect 145010 28590 145012 28642
rect 144956 28588 145012 28590
rect 146076 28028 146132 28084
rect 144284 27746 144340 27748
rect 144284 27694 144286 27746
rect 144286 27694 144338 27746
rect 144338 27694 144340 27746
rect 144284 27692 144340 27694
rect 144956 27692 145012 27748
rect 146076 27132 146132 27188
rect 144396 26962 144452 26964
rect 144396 26910 144398 26962
rect 144398 26910 144450 26962
rect 144450 26910 144452 26962
rect 144396 26908 144452 26910
rect 144956 26908 145012 26964
rect 146076 26236 146132 26292
rect 144396 25282 144452 25284
rect 144396 25230 144398 25282
rect 144398 25230 144450 25282
rect 144450 25230 144452 25282
rect 144396 25228 144452 25230
rect 146076 25394 146132 25396
rect 146076 25342 146078 25394
rect 146078 25342 146130 25394
rect 146130 25342 146132 25394
rect 146076 25340 146132 25342
rect 144956 25228 145012 25284
rect 144284 24610 144340 24612
rect 144284 24558 144286 24610
rect 144286 24558 144338 24610
rect 144338 24558 144340 24610
rect 144284 24556 144340 24558
rect 144956 24556 145012 24612
rect 146076 24444 146132 24500
rect 144396 23714 144452 23716
rect 144396 23662 144398 23714
rect 144398 23662 144450 23714
rect 144450 23662 144452 23714
rect 144396 23660 144452 23662
rect 144956 23660 145012 23716
rect 146076 23660 146132 23716
rect 144284 23042 144340 23044
rect 144284 22990 144286 23042
rect 144286 22990 144338 23042
rect 144338 22990 144340 23042
rect 144284 22988 144340 22990
rect 144956 22988 145012 23044
rect 146076 22652 146132 22708
rect 144396 22146 144452 22148
rect 144396 22094 144398 22146
rect 144398 22094 144450 22146
rect 144450 22094 144452 22146
rect 144396 22092 144452 22094
rect 144956 22092 145012 22148
rect 146076 21756 146132 21812
rect 144284 21474 144340 21476
rect 144284 21422 144286 21474
rect 144286 21422 144338 21474
rect 144338 21422 144340 21474
rect 144284 21420 144340 21422
rect 144956 21420 145012 21476
rect 146076 20860 146132 20916
rect 144396 20578 144452 20580
rect 144396 20526 144398 20578
rect 144398 20526 144450 20578
rect 144450 20526 144452 20578
rect 144396 20524 144452 20526
rect 144956 20524 145012 20580
rect 146076 19964 146132 20020
rect 144396 19010 144452 19012
rect 144396 18958 144398 19010
rect 144398 18958 144450 19010
rect 144450 18958 144452 19010
rect 144396 18956 144452 18958
rect 146076 19122 146132 19124
rect 146076 19070 146078 19122
rect 146078 19070 146130 19122
rect 146130 19070 146132 19122
rect 146076 19068 146132 19070
rect 144956 18956 145012 19012
rect 144284 18338 144340 18340
rect 144284 18286 144286 18338
rect 144286 18286 144338 18338
rect 144338 18286 144340 18338
rect 144284 18284 144340 18286
rect 144956 18284 145012 18340
rect 146076 18172 146132 18228
rect 144396 17442 144452 17444
rect 144396 17390 144398 17442
rect 144398 17390 144450 17442
rect 144450 17390 144452 17442
rect 144396 17388 144452 17390
rect 144956 17388 145012 17444
rect 146076 17388 146132 17444
rect 144284 16882 144340 16884
rect 144284 16830 144286 16882
rect 144286 16830 144338 16882
rect 144338 16830 144340 16882
rect 144284 16828 144340 16830
rect 144956 16882 145012 16884
rect 144956 16830 144958 16882
rect 144958 16830 145010 16882
rect 145010 16830 145012 16882
rect 144956 16828 145012 16830
rect 146076 16380 146132 16436
rect 144396 15874 144452 15876
rect 144396 15822 144398 15874
rect 144398 15822 144450 15874
rect 144450 15822 144452 15874
rect 144396 15820 144452 15822
rect 144956 15820 145012 15876
rect 146076 15484 146132 15540
rect 144284 15260 144340 15316
rect 144956 15314 145012 15316
rect 144956 15262 144958 15314
rect 144958 15262 145010 15314
rect 145010 15262 145012 15314
rect 144956 15260 145012 15262
rect 146076 14588 146132 14644
rect 144396 14306 144452 14308
rect 144396 14254 144398 14306
rect 144398 14254 144450 14306
rect 144450 14254 144452 14306
rect 144396 14252 144452 14254
rect 144956 14252 145012 14308
rect 146076 13692 146132 13748
rect 144284 12796 144340 12852
rect 144396 12908 144452 12964
rect 144956 12962 145012 12964
rect 144956 12910 144958 12962
rect 144958 12910 145010 12962
rect 145010 12910 145012 12962
rect 144956 12908 145012 12910
rect 146076 12850 146132 12852
rect 146076 12798 146078 12850
rect 146078 12798 146130 12850
rect 146130 12798 146132 12850
rect 146076 12796 146132 12798
rect 144284 12066 144340 12068
rect 144284 12014 144286 12066
rect 144286 12014 144338 12066
rect 144338 12014 144340 12066
rect 144284 12012 144340 12014
rect 144620 12236 144676 12292
rect 144284 11116 144340 11172
rect 144396 10780 144452 10836
rect 144284 6578 144340 6580
rect 144284 6526 144286 6578
rect 144286 6526 144338 6578
rect 144338 6526 144340 6578
rect 144284 6524 144340 6526
rect 144956 12012 145012 12068
rect 146076 11900 146132 11956
rect 146076 11116 146132 11172
rect 144956 10780 145012 10836
rect 144956 9938 145012 9940
rect 144956 9886 144958 9938
rect 144958 9886 145010 9938
rect 145010 9886 145012 9938
rect 144956 9884 145012 9886
rect 144956 8930 145012 8932
rect 144956 8878 144958 8930
rect 144958 8878 145010 8930
rect 145010 8878 145012 8930
rect 144956 8876 145012 8878
rect 145068 7756 145124 7812
rect 144956 7420 145012 7476
rect 146300 10108 146356 10164
rect 146860 10108 146916 10164
rect 146300 9714 146356 9716
rect 146300 9662 146302 9714
rect 146302 9662 146354 9714
rect 146354 9662 146356 9714
rect 146300 9660 146356 9662
rect 146972 9660 147028 9716
rect 146972 9212 147028 9268
rect 146300 9154 146356 9156
rect 146300 9102 146302 9154
rect 146302 9102 146354 9154
rect 146354 9102 146356 9154
rect 146300 9100 146356 9102
rect 146860 9100 146916 9156
rect 146860 8428 146916 8484
rect 146300 8146 146356 8148
rect 146300 8094 146302 8146
rect 146302 8094 146354 8146
rect 146354 8094 146356 8146
rect 146300 8092 146356 8094
rect 146972 8092 147028 8148
rect 145180 7532 145236 7588
rect 146188 7586 146244 7588
rect 146188 7534 146190 7586
rect 146190 7534 146242 7586
rect 146242 7534 146244 7586
rect 146188 7532 146244 7534
rect 144732 6636 144788 6692
rect 145180 6524 145236 6580
rect 144956 6188 145012 6244
rect 144620 4956 144676 5012
rect 144172 3442 144228 3444
rect 144172 3390 144174 3442
rect 144174 3390 144226 3442
rect 144226 3390 144228 3442
rect 144172 3388 144228 3390
rect 143948 2492 144004 2548
rect 144956 4226 145012 4228
rect 144956 4174 144958 4226
rect 144958 4174 145010 4226
rect 145010 4174 145012 4226
rect 144956 4172 145012 4174
rect 145068 3442 145124 3444
rect 145068 3390 145070 3442
rect 145070 3390 145122 3442
rect 145122 3390 145124 3442
rect 145068 3388 145124 3390
rect 145180 2940 145236 2996
rect 145964 5740 146020 5796
rect 146860 7586 146916 7588
rect 146860 7534 146862 7586
rect 146862 7534 146914 7586
rect 146914 7534 146916 7586
rect 146860 7532 146916 7534
rect 147084 7644 147140 7700
rect 147868 34636 147924 34692
rect 146972 7420 147028 7476
rect 146300 6578 146356 6580
rect 146300 6526 146302 6578
rect 146302 6526 146354 6578
rect 146354 6526 146356 6578
rect 146300 6524 146356 6526
rect 146972 6578 147028 6580
rect 146972 6526 146974 6578
rect 146974 6526 147026 6578
rect 147026 6526 147028 6578
rect 146972 6524 147028 6526
rect 146860 5794 146916 5796
rect 146860 5742 146862 5794
rect 146862 5742 146914 5794
rect 146914 5742 146916 5794
rect 146860 5740 146916 5742
rect 146300 5628 146356 5684
rect 147308 5628 147364 5684
rect 146860 4956 146916 5012
rect 146300 4844 146356 4900
rect 147420 4898 147476 4900
rect 147420 4846 147422 4898
rect 147422 4846 147474 4898
rect 147474 4846 147476 4898
rect 147420 4844 147476 4846
rect 146300 3836 146356 3892
rect 146860 3836 146916 3892
rect 148492 34522 148548 34524
rect 148492 34470 148494 34522
rect 148494 34470 148546 34522
rect 148546 34470 148548 34522
rect 148492 34468 148548 34470
rect 148596 34522 148652 34524
rect 148596 34470 148598 34522
rect 148598 34470 148650 34522
rect 148650 34470 148652 34522
rect 148596 34468 148652 34470
rect 148700 34522 148756 34524
rect 148700 34470 148702 34522
rect 148702 34470 148754 34522
rect 148754 34470 148756 34522
rect 148700 34468 148756 34470
rect 148492 32954 148548 32956
rect 148492 32902 148494 32954
rect 148494 32902 148546 32954
rect 148546 32902 148548 32954
rect 148492 32900 148548 32902
rect 148596 32954 148652 32956
rect 148596 32902 148598 32954
rect 148598 32902 148650 32954
rect 148650 32902 148652 32954
rect 148596 32900 148652 32902
rect 148700 32954 148756 32956
rect 148700 32902 148702 32954
rect 148702 32902 148754 32954
rect 148754 32902 148756 32954
rect 148700 32900 148756 32902
rect 148492 31386 148548 31388
rect 148492 31334 148494 31386
rect 148494 31334 148546 31386
rect 148546 31334 148548 31386
rect 148492 31332 148548 31334
rect 148596 31386 148652 31388
rect 148596 31334 148598 31386
rect 148598 31334 148650 31386
rect 148650 31334 148652 31386
rect 148596 31332 148652 31334
rect 148700 31386 148756 31388
rect 148700 31334 148702 31386
rect 148702 31334 148754 31386
rect 148754 31334 148756 31386
rect 148700 31332 148756 31334
rect 148492 29818 148548 29820
rect 148492 29766 148494 29818
rect 148494 29766 148546 29818
rect 148546 29766 148548 29818
rect 148492 29764 148548 29766
rect 148596 29818 148652 29820
rect 148596 29766 148598 29818
rect 148598 29766 148650 29818
rect 148650 29766 148652 29818
rect 148596 29764 148652 29766
rect 148700 29818 148756 29820
rect 148700 29766 148702 29818
rect 148702 29766 148754 29818
rect 148754 29766 148756 29818
rect 148700 29764 148756 29766
rect 148492 28250 148548 28252
rect 148492 28198 148494 28250
rect 148494 28198 148546 28250
rect 148546 28198 148548 28250
rect 148492 28196 148548 28198
rect 148596 28250 148652 28252
rect 148596 28198 148598 28250
rect 148598 28198 148650 28250
rect 148650 28198 148652 28250
rect 148596 28196 148652 28198
rect 148700 28250 148756 28252
rect 148700 28198 148702 28250
rect 148702 28198 148754 28250
rect 148754 28198 148756 28250
rect 148700 28196 148756 28198
rect 148492 26682 148548 26684
rect 148492 26630 148494 26682
rect 148494 26630 148546 26682
rect 148546 26630 148548 26682
rect 148492 26628 148548 26630
rect 148596 26682 148652 26684
rect 148596 26630 148598 26682
rect 148598 26630 148650 26682
rect 148650 26630 148652 26682
rect 148596 26628 148652 26630
rect 148700 26682 148756 26684
rect 148700 26630 148702 26682
rect 148702 26630 148754 26682
rect 148754 26630 148756 26682
rect 148700 26628 148756 26630
rect 148492 25114 148548 25116
rect 148492 25062 148494 25114
rect 148494 25062 148546 25114
rect 148546 25062 148548 25114
rect 148492 25060 148548 25062
rect 148596 25114 148652 25116
rect 148596 25062 148598 25114
rect 148598 25062 148650 25114
rect 148650 25062 148652 25114
rect 148596 25060 148652 25062
rect 148700 25114 148756 25116
rect 148700 25062 148702 25114
rect 148702 25062 148754 25114
rect 148754 25062 148756 25114
rect 148700 25060 148756 25062
rect 148492 23546 148548 23548
rect 148492 23494 148494 23546
rect 148494 23494 148546 23546
rect 148546 23494 148548 23546
rect 148492 23492 148548 23494
rect 148596 23546 148652 23548
rect 148596 23494 148598 23546
rect 148598 23494 148650 23546
rect 148650 23494 148652 23546
rect 148596 23492 148652 23494
rect 148700 23546 148756 23548
rect 148700 23494 148702 23546
rect 148702 23494 148754 23546
rect 148754 23494 148756 23546
rect 148700 23492 148756 23494
rect 148492 21978 148548 21980
rect 148492 21926 148494 21978
rect 148494 21926 148546 21978
rect 148546 21926 148548 21978
rect 148492 21924 148548 21926
rect 148596 21978 148652 21980
rect 148596 21926 148598 21978
rect 148598 21926 148650 21978
rect 148650 21926 148652 21978
rect 148596 21924 148652 21926
rect 148700 21978 148756 21980
rect 148700 21926 148702 21978
rect 148702 21926 148754 21978
rect 148754 21926 148756 21978
rect 148700 21924 148756 21926
rect 148492 20410 148548 20412
rect 148492 20358 148494 20410
rect 148494 20358 148546 20410
rect 148546 20358 148548 20410
rect 148492 20356 148548 20358
rect 148596 20410 148652 20412
rect 148596 20358 148598 20410
rect 148598 20358 148650 20410
rect 148650 20358 148652 20410
rect 148596 20356 148652 20358
rect 148700 20410 148756 20412
rect 148700 20358 148702 20410
rect 148702 20358 148754 20410
rect 148754 20358 148756 20410
rect 148700 20356 148756 20358
rect 148492 18842 148548 18844
rect 148492 18790 148494 18842
rect 148494 18790 148546 18842
rect 148546 18790 148548 18842
rect 148492 18788 148548 18790
rect 148596 18842 148652 18844
rect 148596 18790 148598 18842
rect 148598 18790 148650 18842
rect 148650 18790 148652 18842
rect 148596 18788 148652 18790
rect 148700 18842 148756 18844
rect 148700 18790 148702 18842
rect 148702 18790 148754 18842
rect 148754 18790 148756 18842
rect 148700 18788 148756 18790
rect 148492 17274 148548 17276
rect 148492 17222 148494 17274
rect 148494 17222 148546 17274
rect 148546 17222 148548 17274
rect 148492 17220 148548 17222
rect 148596 17274 148652 17276
rect 148596 17222 148598 17274
rect 148598 17222 148650 17274
rect 148650 17222 148652 17274
rect 148596 17220 148652 17222
rect 148700 17274 148756 17276
rect 148700 17222 148702 17274
rect 148702 17222 148754 17274
rect 148754 17222 148756 17274
rect 148700 17220 148756 17222
rect 148492 15706 148548 15708
rect 148492 15654 148494 15706
rect 148494 15654 148546 15706
rect 148546 15654 148548 15706
rect 148492 15652 148548 15654
rect 148596 15706 148652 15708
rect 148596 15654 148598 15706
rect 148598 15654 148650 15706
rect 148650 15654 148652 15706
rect 148596 15652 148652 15654
rect 148700 15706 148756 15708
rect 148700 15654 148702 15706
rect 148702 15654 148754 15706
rect 148754 15654 148756 15706
rect 148700 15652 148756 15654
rect 148492 14138 148548 14140
rect 148492 14086 148494 14138
rect 148494 14086 148546 14138
rect 148546 14086 148548 14138
rect 148492 14084 148548 14086
rect 148596 14138 148652 14140
rect 148596 14086 148598 14138
rect 148598 14086 148650 14138
rect 148650 14086 148652 14138
rect 148596 14084 148652 14086
rect 148700 14138 148756 14140
rect 148700 14086 148702 14138
rect 148702 14086 148754 14138
rect 148754 14086 148756 14138
rect 148700 14084 148756 14086
rect 148492 12570 148548 12572
rect 148492 12518 148494 12570
rect 148494 12518 148546 12570
rect 148546 12518 148548 12570
rect 148492 12516 148548 12518
rect 148596 12570 148652 12572
rect 148596 12518 148598 12570
rect 148598 12518 148650 12570
rect 148650 12518 148652 12570
rect 148596 12516 148652 12518
rect 148700 12570 148756 12572
rect 148700 12518 148702 12570
rect 148702 12518 148754 12570
rect 148754 12518 148756 12570
rect 148700 12516 148756 12518
rect 148492 11002 148548 11004
rect 148492 10950 148494 11002
rect 148494 10950 148546 11002
rect 148546 10950 148548 11002
rect 148492 10948 148548 10950
rect 148596 11002 148652 11004
rect 148596 10950 148598 11002
rect 148598 10950 148650 11002
rect 148650 10950 148652 11002
rect 148596 10948 148652 10950
rect 148700 11002 148756 11004
rect 148700 10950 148702 11002
rect 148702 10950 148754 11002
rect 148754 10950 148756 11002
rect 148700 10948 148756 10950
rect 148492 9434 148548 9436
rect 148492 9382 148494 9434
rect 148494 9382 148546 9434
rect 148546 9382 148548 9434
rect 148492 9380 148548 9382
rect 148596 9434 148652 9436
rect 148596 9382 148598 9434
rect 148598 9382 148650 9434
rect 148650 9382 148652 9434
rect 148596 9380 148652 9382
rect 148700 9434 148756 9436
rect 148700 9382 148702 9434
rect 148702 9382 148754 9434
rect 148754 9382 148756 9434
rect 148700 9380 148756 9382
rect 148492 7866 148548 7868
rect 148492 7814 148494 7866
rect 148494 7814 148546 7866
rect 148546 7814 148548 7866
rect 148492 7812 148548 7814
rect 148596 7866 148652 7868
rect 148596 7814 148598 7866
rect 148598 7814 148650 7866
rect 148650 7814 148652 7866
rect 148596 7812 148652 7814
rect 148700 7866 148756 7868
rect 148700 7814 148702 7866
rect 148702 7814 148754 7866
rect 148754 7814 148756 7866
rect 148700 7812 148756 7814
rect 148492 6298 148548 6300
rect 148492 6246 148494 6298
rect 148494 6246 148546 6298
rect 148546 6246 148548 6298
rect 148492 6244 148548 6246
rect 148596 6298 148652 6300
rect 148596 6246 148598 6298
rect 148598 6246 148650 6298
rect 148650 6246 148652 6298
rect 148596 6244 148652 6246
rect 148700 6298 148756 6300
rect 148700 6246 148702 6298
rect 148702 6246 148754 6298
rect 148754 6246 148756 6298
rect 148700 6244 148756 6246
rect 148492 4730 148548 4732
rect 148492 4678 148494 4730
rect 148494 4678 148546 4730
rect 148546 4678 148548 4730
rect 148492 4676 148548 4678
rect 148596 4730 148652 4732
rect 148596 4678 148598 4730
rect 148598 4678 148650 4730
rect 148650 4678 148652 4730
rect 148596 4676 148652 4678
rect 148700 4730 148756 4732
rect 148700 4678 148702 4730
rect 148702 4678 148754 4730
rect 148754 4678 148756 4730
rect 148700 4676 148756 4678
rect 147868 3276 147924 3332
rect 148492 3162 148548 3164
rect 148492 3110 148494 3162
rect 148494 3110 148546 3162
rect 148546 3110 148548 3162
rect 148492 3108 148548 3110
rect 148596 3162 148652 3164
rect 148596 3110 148598 3162
rect 148598 3110 148650 3162
rect 148650 3110 148652 3162
rect 148596 3108 148652 3110
rect 148700 3162 148756 3164
rect 148700 3110 148702 3162
rect 148702 3110 148754 3162
rect 148754 3110 148756 3162
rect 148700 3108 148756 3110
rect 146076 2044 146132 2100
rect 145964 1148 146020 1204
<< metal3 >>
rect 149200 38836 150000 38864
rect 147634 38780 147644 38836
rect 147700 38780 150000 38836
rect 149200 38752 150000 38780
rect 149200 37940 150000 37968
rect 144498 37884 144508 37940
rect 144564 37884 150000 37940
rect 149200 37856 150000 37884
rect 149200 37044 150000 37072
rect 147746 36988 147756 37044
rect 147812 36988 150000 37044
rect 149200 36960 150000 36988
rect 19612 36820 19622 36876
rect 19678 36820 19726 36876
rect 19782 36820 19830 36876
rect 19886 36820 19896 36876
rect 56432 36820 56442 36876
rect 56498 36820 56546 36876
rect 56602 36820 56650 36876
rect 56706 36820 56716 36876
rect 93252 36820 93262 36876
rect 93318 36820 93366 36876
rect 93422 36820 93470 36876
rect 93526 36820 93536 36876
rect 130072 36820 130082 36876
rect 130138 36820 130186 36876
rect 130242 36820 130290 36876
rect 130346 36820 130356 36876
rect 144162 36316 144172 36372
rect 144228 36316 144844 36372
rect 144900 36316 144910 36372
rect 139010 36204 139020 36260
rect 139076 36204 142156 36260
rect 142212 36204 143052 36260
rect 143108 36204 143118 36260
rect 145954 36204 145964 36260
rect 146020 36204 148932 36260
rect 148876 36148 148932 36204
rect 149200 36148 150000 36176
rect 148876 36092 150000 36148
rect 38022 36036 38032 36092
rect 38088 36036 38136 36092
rect 38192 36036 38240 36092
rect 38296 36036 38306 36092
rect 74842 36036 74852 36092
rect 74908 36036 74956 36092
rect 75012 36036 75060 36092
rect 75116 36036 75126 36092
rect 111662 36036 111672 36092
rect 111728 36036 111776 36092
rect 111832 36036 111880 36092
rect 111936 36036 111946 36092
rect 148482 36036 148492 36092
rect 148548 36036 148596 36092
rect 148652 36036 148700 36092
rect 148756 36036 148766 36092
rect 149200 36064 150000 36092
rect 142146 35532 142156 35588
rect 142212 35532 144284 35588
rect 144340 35532 144956 35588
rect 145012 35532 145022 35588
rect 19612 35252 19622 35308
rect 19678 35252 19726 35308
rect 19782 35252 19830 35308
rect 19886 35252 19896 35308
rect 56432 35252 56442 35308
rect 56498 35252 56546 35308
rect 56602 35252 56650 35308
rect 56706 35252 56716 35308
rect 93252 35252 93262 35308
rect 93318 35252 93366 35308
rect 93422 35252 93470 35308
rect 93526 35252 93536 35308
rect 130072 35252 130082 35308
rect 130138 35252 130186 35308
rect 130242 35252 130290 35308
rect 130346 35252 130356 35308
rect 149200 35252 150000 35280
rect 146066 35196 146076 35252
rect 146132 35196 150000 35252
rect 149200 35168 150000 35196
rect 141250 34636 141260 34692
rect 141316 34636 144396 34692
rect 144452 34636 144956 34692
rect 145012 34636 145022 34692
rect 146626 34636 146636 34692
rect 146692 34636 147868 34692
rect 147924 34636 147934 34692
rect 38022 34468 38032 34524
rect 38088 34468 38136 34524
rect 38192 34468 38240 34524
rect 38296 34468 38306 34524
rect 74842 34468 74852 34524
rect 74908 34468 74956 34524
rect 75012 34468 75060 34524
rect 75116 34468 75126 34524
rect 111662 34468 111672 34524
rect 111728 34468 111776 34524
rect 111832 34468 111880 34524
rect 111936 34468 111946 34524
rect 148482 34468 148492 34524
rect 148548 34468 148596 34524
rect 148652 34468 148700 34524
rect 148756 34468 148766 34524
rect 149200 34356 150000 34384
rect 146066 34300 146076 34356
rect 146132 34300 150000 34356
rect 149200 34272 150000 34300
rect 137330 33964 137340 34020
rect 137396 33964 144284 34020
rect 144340 33964 144956 34020
rect 145012 33964 145022 34020
rect 19612 33684 19622 33740
rect 19678 33684 19726 33740
rect 19782 33684 19830 33740
rect 19886 33684 19896 33740
rect 56432 33684 56442 33740
rect 56498 33684 56546 33740
rect 56602 33684 56650 33740
rect 56706 33684 56716 33740
rect 93252 33684 93262 33740
rect 93318 33684 93366 33740
rect 93422 33684 93470 33740
rect 93526 33684 93536 33740
rect 130072 33684 130082 33740
rect 130138 33684 130186 33740
rect 130242 33684 130290 33740
rect 130346 33684 130356 33740
rect 149200 33460 150000 33488
rect 146066 33404 146076 33460
rect 146132 33404 150000 33460
rect 149200 33376 150000 33404
rect 134754 33068 134764 33124
rect 134820 33068 144396 33124
rect 144452 33068 144956 33124
rect 145012 33068 145022 33124
rect 38022 32900 38032 32956
rect 38088 32900 38136 32956
rect 38192 32900 38240 32956
rect 38296 32900 38306 32956
rect 74842 32900 74852 32956
rect 74908 32900 74956 32956
rect 75012 32900 75060 32956
rect 75116 32900 75126 32956
rect 111662 32900 111672 32956
rect 111728 32900 111776 32956
rect 111832 32900 111880 32956
rect 111936 32900 111946 32956
rect 148482 32900 148492 32956
rect 148548 32900 148596 32956
rect 148652 32900 148700 32956
rect 148756 32900 148766 32956
rect 149200 32564 150000 32592
rect 146066 32508 146076 32564
rect 146132 32508 150000 32564
rect 149200 32480 150000 32508
rect 19612 32116 19622 32172
rect 19678 32116 19726 32172
rect 19782 32116 19830 32172
rect 19886 32116 19896 32172
rect 56432 32116 56442 32172
rect 56498 32116 56546 32172
rect 56602 32116 56650 32172
rect 56706 32116 56716 32172
rect 93252 32116 93262 32172
rect 93318 32116 93366 32172
rect 93422 32116 93470 32172
rect 93526 32116 93536 32172
rect 130072 32116 130082 32172
rect 130138 32116 130186 32172
rect 130242 32116 130290 32172
rect 130346 32116 130356 32172
rect 149200 31668 150000 31696
rect 146066 31612 146076 31668
rect 146132 31612 150000 31668
rect 149200 31584 150000 31612
rect 133298 31500 133308 31556
rect 133364 31500 144396 31556
rect 144452 31500 144956 31556
rect 145012 31500 145022 31556
rect 38022 31332 38032 31388
rect 38088 31332 38136 31388
rect 38192 31332 38240 31388
rect 38296 31332 38306 31388
rect 74842 31332 74852 31388
rect 74908 31332 74956 31388
rect 75012 31332 75060 31388
rect 75116 31332 75126 31388
rect 111662 31332 111672 31388
rect 111728 31332 111776 31388
rect 111832 31332 111880 31388
rect 111936 31332 111946 31388
rect 148482 31332 148492 31388
rect 148548 31332 148596 31388
rect 148652 31332 148700 31388
rect 148756 31332 148766 31388
rect 131394 30828 131404 30884
rect 131460 30828 144284 30884
rect 144340 30828 144956 30884
rect 145012 30828 145022 30884
rect 149200 30772 150000 30800
rect 146066 30716 146076 30772
rect 146132 30716 150000 30772
rect 149200 30688 150000 30716
rect 19612 30548 19622 30604
rect 19678 30548 19726 30604
rect 19782 30548 19830 30604
rect 19886 30548 19896 30604
rect 56432 30548 56442 30604
rect 56498 30548 56546 30604
rect 56602 30548 56650 30604
rect 56706 30548 56716 30604
rect 93252 30548 93262 30604
rect 93318 30548 93366 30604
rect 93422 30548 93470 30604
rect 93526 30548 93536 30604
rect 130072 30548 130082 30604
rect 130138 30548 130186 30604
rect 130242 30548 130290 30604
rect 130346 30548 130356 30604
rect 138562 29932 138572 29988
rect 138628 29932 144396 29988
rect 144452 29932 144956 29988
rect 145012 29932 145022 29988
rect 146066 29932 146076 29988
rect 146132 29932 148932 29988
rect 148876 29876 148932 29932
rect 149200 29876 150000 29904
rect 148876 29820 150000 29876
rect 38022 29764 38032 29820
rect 38088 29764 38136 29820
rect 38192 29764 38240 29820
rect 38296 29764 38306 29820
rect 74842 29764 74852 29820
rect 74908 29764 74956 29820
rect 75012 29764 75060 29820
rect 75116 29764 75126 29820
rect 111662 29764 111672 29820
rect 111728 29764 111776 29820
rect 111832 29764 111880 29820
rect 111936 29764 111946 29820
rect 148482 29764 148492 29820
rect 148548 29764 148596 29820
rect 148652 29764 148700 29820
rect 148756 29764 148766 29820
rect 149200 29792 150000 29820
rect 127922 29260 127932 29316
rect 127988 29260 144284 29316
rect 144340 29260 144956 29316
rect 145012 29260 145022 29316
rect 19612 28980 19622 29036
rect 19678 28980 19726 29036
rect 19782 28980 19830 29036
rect 19886 28980 19896 29036
rect 56432 28980 56442 29036
rect 56498 28980 56546 29036
rect 56602 28980 56650 29036
rect 56706 28980 56716 29036
rect 93252 28980 93262 29036
rect 93318 28980 93366 29036
rect 93422 28980 93470 29036
rect 93526 28980 93536 29036
rect 130072 28980 130082 29036
rect 130138 28980 130186 29036
rect 130242 28980 130290 29036
rect 130346 28980 130356 29036
rect 149200 28980 150000 29008
rect 146066 28924 146076 28980
rect 146132 28924 150000 28980
rect 149200 28896 150000 28924
rect 141026 28588 141036 28644
rect 141092 28588 144396 28644
rect 144452 28588 144956 28644
rect 145012 28588 145022 28644
rect 38022 28196 38032 28252
rect 38088 28196 38136 28252
rect 38192 28196 38240 28252
rect 38296 28196 38306 28252
rect 74842 28196 74852 28252
rect 74908 28196 74956 28252
rect 75012 28196 75060 28252
rect 75116 28196 75126 28252
rect 111662 28196 111672 28252
rect 111728 28196 111776 28252
rect 111832 28196 111880 28252
rect 111936 28196 111946 28252
rect 148482 28196 148492 28252
rect 148548 28196 148596 28252
rect 148652 28196 148700 28252
rect 148756 28196 148766 28252
rect 149200 28084 150000 28112
rect 146066 28028 146076 28084
rect 146132 28028 150000 28084
rect 149200 28000 150000 28028
rect 124898 27692 124908 27748
rect 124964 27692 144284 27748
rect 144340 27692 144956 27748
rect 145012 27692 145022 27748
rect 19612 27412 19622 27468
rect 19678 27412 19726 27468
rect 19782 27412 19830 27468
rect 19886 27412 19896 27468
rect 56432 27412 56442 27468
rect 56498 27412 56546 27468
rect 56602 27412 56650 27468
rect 56706 27412 56716 27468
rect 93252 27412 93262 27468
rect 93318 27412 93366 27468
rect 93422 27412 93470 27468
rect 93526 27412 93536 27468
rect 130072 27412 130082 27468
rect 130138 27412 130186 27468
rect 130242 27412 130290 27468
rect 130346 27412 130356 27468
rect 149200 27188 150000 27216
rect 146066 27132 146076 27188
rect 146132 27132 150000 27188
rect 149200 27104 150000 27132
rect 124114 26908 124124 26964
rect 124180 26908 144396 26964
rect 144452 26908 144956 26964
rect 145012 26908 145022 26964
rect 38022 26628 38032 26684
rect 38088 26628 38136 26684
rect 38192 26628 38240 26684
rect 38296 26628 38306 26684
rect 74842 26628 74852 26684
rect 74908 26628 74956 26684
rect 75012 26628 75060 26684
rect 75116 26628 75126 26684
rect 111662 26628 111672 26684
rect 111728 26628 111776 26684
rect 111832 26628 111880 26684
rect 111936 26628 111946 26684
rect 148482 26628 148492 26684
rect 148548 26628 148596 26684
rect 148652 26628 148700 26684
rect 148756 26628 148766 26684
rect 149200 26292 150000 26320
rect 146066 26236 146076 26292
rect 146132 26236 150000 26292
rect 149200 26208 150000 26236
rect 19612 25844 19622 25900
rect 19678 25844 19726 25900
rect 19782 25844 19830 25900
rect 19886 25844 19896 25900
rect 56432 25844 56442 25900
rect 56498 25844 56546 25900
rect 56602 25844 56650 25900
rect 56706 25844 56716 25900
rect 93252 25844 93262 25900
rect 93318 25844 93366 25900
rect 93422 25844 93470 25900
rect 93526 25844 93536 25900
rect 130072 25844 130082 25900
rect 130138 25844 130186 25900
rect 130242 25844 130290 25900
rect 130346 25844 130356 25900
rect 149200 25396 150000 25424
rect 146066 25340 146076 25396
rect 146132 25340 150000 25396
rect 149200 25312 150000 25340
rect 122220 25228 144396 25284
rect 144452 25228 144956 25284
rect 145012 25228 145022 25284
rect 122220 25172 122276 25228
rect 120082 25116 120092 25172
rect 120148 25116 122276 25172
rect 38022 25060 38032 25116
rect 38088 25060 38136 25116
rect 38192 25060 38240 25116
rect 38296 25060 38306 25116
rect 74842 25060 74852 25116
rect 74908 25060 74956 25116
rect 75012 25060 75060 25116
rect 75116 25060 75126 25116
rect 111662 25060 111672 25116
rect 111728 25060 111776 25116
rect 111832 25060 111880 25116
rect 111936 25060 111946 25116
rect 148482 25060 148492 25116
rect 148548 25060 148596 25116
rect 148652 25060 148700 25116
rect 148756 25060 148766 25116
rect 119186 24556 119196 24612
rect 119252 24556 144284 24612
rect 144340 24556 144956 24612
rect 145012 24556 145022 24612
rect 149200 24500 150000 24528
rect 146066 24444 146076 24500
rect 146132 24444 150000 24500
rect 149200 24416 150000 24444
rect 19612 24276 19622 24332
rect 19678 24276 19726 24332
rect 19782 24276 19830 24332
rect 19886 24276 19896 24332
rect 56432 24276 56442 24332
rect 56498 24276 56546 24332
rect 56602 24276 56650 24332
rect 56706 24276 56716 24332
rect 93252 24276 93262 24332
rect 93318 24276 93366 24332
rect 93422 24276 93470 24332
rect 93526 24276 93536 24332
rect 130072 24276 130082 24332
rect 130138 24276 130186 24332
rect 130242 24276 130290 24332
rect 130346 24276 130356 24332
rect 121762 23660 121772 23716
rect 121828 23660 144396 23716
rect 144452 23660 144956 23716
rect 145012 23660 145022 23716
rect 146066 23660 146076 23716
rect 146132 23660 148932 23716
rect 148876 23604 148932 23660
rect 149200 23604 150000 23632
rect 148876 23548 150000 23604
rect 38022 23492 38032 23548
rect 38088 23492 38136 23548
rect 38192 23492 38240 23548
rect 38296 23492 38306 23548
rect 74842 23492 74852 23548
rect 74908 23492 74956 23548
rect 75012 23492 75060 23548
rect 75116 23492 75126 23548
rect 111662 23492 111672 23548
rect 111728 23492 111776 23548
rect 111832 23492 111880 23548
rect 111936 23492 111946 23548
rect 148482 23492 148492 23548
rect 148548 23492 148596 23548
rect 148652 23492 148700 23548
rect 148756 23492 148766 23548
rect 149200 23520 150000 23548
rect 139458 22988 139468 23044
rect 139524 22988 144284 23044
rect 144340 22988 144956 23044
rect 145012 22988 145022 23044
rect 126018 22876 126028 22932
rect 126084 22876 141036 22932
rect 141092 22876 141102 22932
rect 19612 22708 19622 22764
rect 19678 22708 19726 22764
rect 19782 22708 19830 22764
rect 19886 22708 19896 22764
rect 56432 22708 56442 22764
rect 56498 22708 56546 22764
rect 56602 22708 56650 22764
rect 56706 22708 56716 22764
rect 93252 22708 93262 22764
rect 93318 22708 93366 22764
rect 93422 22708 93470 22764
rect 93526 22708 93536 22764
rect 130072 22708 130082 22764
rect 130138 22708 130186 22764
rect 130242 22708 130290 22764
rect 130346 22708 130356 22764
rect 149200 22708 150000 22736
rect 146066 22652 146076 22708
rect 146132 22652 150000 22708
rect 149200 22624 150000 22652
rect 113474 22092 113484 22148
rect 113540 22092 144396 22148
rect 144452 22092 144956 22148
rect 145012 22092 145022 22148
rect 38022 21924 38032 21980
rect 38088 21924 38136 21980
rect 38192 21924 38240 21980
rect 38296 21924 38306 21980
rect 74842 21924 74852 21980
rect 74908 21924 74956 21980
rect 75012 21924 75060 21980
rect 75116 21924 75126 21980
rect 111662 21924 111672 21980
rect 111728 21924 111776 21980
rect 111832 21924 111880 21980
rect 111936 21924 111946 21980
rect 148482 21924 148492 21980
rect 148548 21924 148596 21980
rect 148652 21924 148700 21980
rect 148756 21924 148766 21980
rect 149200 21812 150000 21840
rect 146066 21756 146076 21812
rect 146132 21756 150000 21812
rect 149200 21728 150000 21756
rect 143490 21420 143500 21476
rect 143556 21420 144284 21476
rect 144340 21420 144956 21476
rect 145012 21420 145022 21476
rect 19612 21140 19622 21196
rect 19678 21140 19726 21196
rect 19782 21140 19830 21196
rect 19886 21140 19896 21196
rect 56432 21140 56442 21196
rect 56498 21140 56546 21196
rect 56602 21140 56650 21196
rect 56706 21140 56716 21196
rect 93252 21140 93262 21196
rect 93318 21140 93366 21196
rect 93422 21140 93470 21196
rect 93526 21140 93536 21196
rect 130072 21140 130082 21196
rect 130138 21140 130186 21196
rect 130242 21140 130290 21196
rect 130346 21140 130356 21196
rect 149200 20916 150000 20944
rect 146066 20860 146076 20916
rect 146132 20860 150000 20916
rect 149200 20832 150000 20860
rect 114258 20524 114268 20580
rect 114324 20524 144396 20580
rect 144452 20524 144956 20580
rect 145012 20524 145022 20580
rect 38022 20356 38032 20412
rect 38088 20356 38136 20412
rect 38192 20356 38240 20412
rect 38296 20356 38306 20412
rect 74842 20356 74852 20412
rect 74908 20356 74956 20412
rect 75012 20356 75060 20412
rect 75116 20356 75126 20412
rect 111662 20356 111672 20412
rect 111728 20356 111776 20412
rect 111832 20356 111880 20412
rect 111936 20356 111946 20412
rect 148482 20356 148492 20412
rect 148548 20356 148596 20412
rect 148652 20356 148700 20412
rect 148756 20356 148766 20412
rect 149200 20020 150000 20048
rect 146066 19964 146076 20020
rect 146132 19964 150000 20020
rect 149200 19936 150000 19964
rect 19612 19572 19622 19628
rect 19678 19572 19726 19628
rect 19782 19572 19830 19628
rect 19886 19572 19896 19628
rect 56432 19572 56442 19628
rect 56498 19572 56546 19628
rect 56602 19572 56650 19628
rect 56706 19572 56716 19628
rect 93252 19572 93262 19628
rect 93318 19572 93366 19628
rect 93422 19572 93470 19628
rect 93526 19572 93536 19628
rect 130072 19572 130082 19628
rect 130138 19572 130186 19628
rect 130242 19572 130290 19628
rect 130346 19572 130356 19628
rect 149200 19124 150000 19152
rect 146066 19068 146076 19124
rect 146132 19068 150000 19124
rect 149200 19040 150000 19068
rect 143938 18956 143948 19012
rect 144004 18956 144396 19012
rect 144452 18956 144956 19012
rect 145012 18956 145022 19012
rect 38022 18788 38032 18844
rect 38088 18788 38136 18844
rect 38192 18788 38240 18844
rect 38296 18788 38306 18844
rect 74842 18788 74852 18844
rect 74908 18788 74956 18844
rect 75012 18788 75060 18844
rect 75116 18788 75126 18844
rect 111662 18788 111672 18844
rect 111728 18788 111776 18844
rect 111832 18788 111880 18844
rect 111936 18788 111946 18844
rect 148482 18788 148492 18844
rect 148548 18788 148596 18844
rect 148652 18788 148700 18844
rect 148756 18788 148766 18844
rect 111570 18620 111580 18676
rect 111636 18620 114268 18676
rect 114324 18620 114334 18676
rect 115826 18284 115836 18340
rect 115892 18284 144284 18340
rect 144340 18284 144956 18340
rect 145012 18284 145022 18340
rect 149200 18228 150000 18256
rect 146066 18172 146076 18228
rect 146132 18172 150000 18228
rect 149200 18144 150000 18172
rect 19612 18004 19622 18060
rect 19678 18004 19726 18060
rect 19782 18004 19830 18060
rect 19886 18004 19896 18060
rect 56432 18004 56442 18060
rect 56498 18004 56546 18060
rect 56602 18004 56650 18060
rect 56706 18004 56716 18060
rect 93252 18004 93262 18060
rect 93318 18004 93366 18060
rect 93422 18004 93470 18060
rect 93526 18004 93536 18060
rect 130072 18004 130082 18060
rect 130138 18004 130186 18060
rect 130242 18004 130290 18060
rect 130346 18004 130356 18060
rect 106642 17388 106652 17444
rect 106708 17388 144396 17444
rect 144452 17388 144956 17444
rect 145012 17388 145022 17444
rect 146066 17388 146076 17444
rect 146132 17388 148932 17444
rect 148876 17332 148932 17388
rect 149200 17332 150000 17360
rect 148876 17276 150000 17332
rect 38022 17220 38032 17276
rect 38088 17220 38136 17276
rect 38192 17220 38240 17276
rect 38296 17220 38306 17276
rect 74842 17220 74852 17276
rect 74908 17220 74956 17276
rect 75012 17220 75060 17276
rect 75116 17220 75126 17276
rect 111662 17220 111672 17276
rect 111728 17220 111776 17276
rect 111832 17220 111880 17276
rect 111936 17220 111946 17276
rect 148482 17220 148492 17276
rect 148548 17220 148596 17276
rect 148652 17220 148700 17276
rect 148756 17220 148766 17276
rect 149200 17248 150000 17276
rect 104514 16828 104524 16884
rect 104580 16828 144284 16884
rect 144340 16828 144956 16884
rect 145012 16828 145022 16884
rect 19612 16436 19622 16492
rect 19678 16436 19726 16492
rect 19782 16436 19830 16492
rect 19886 16436 19896 16492
rect 56432 16436 56442 16492
rect 56498 16436 56546 16492
rect 56602 16436 56650 16492
rect 56706 16436 56716 16492
rect 93252 16436 93262 16492
rect 93318 16436 93366 16492
rect 93422 16436 93470 16492
rect 93526 16436 93536 16492
rect 130072 16436 130082 16492
rect 130138 16436 130186 16492
rect 130242 16436 130290 16492
rect 130346 16436 130356 16492
rect 149200 16436 150000 16464
rect 146066 16380 146076 16436
rect 146132 16380 150000 16436
rect 149200 16352 150000 16380
rect 103618 15820 103628 15876
rect 103684 15820 144396 15876
rect 144452 15820 144956 15876
rect 145012 15820 145022 15876
rect 38022 15652 38032 15708
rect 38088 15652 38136 15708
rect 38192 15652 38240 15708
rect 38296 15652 38306 15708
rect 74842 15652 74852 15708
rect 74908 15652 74956 15708
rect 75012 15652 75060 15708
rect 75116 15652 75126 15708
rect 111662 15652 111672 15708
rect 111728 15652 111776 15708
rect 111832 15652 111880 15708
rect 111936 15652 111946 15708
rect 148482 15652 148492 15708
rect 148548 15652 148596 15708
rect 148652 15652 148700 15708
rect 148756 15652 148766 15708
rect 149200 15540 150000 15568
rect 146066 15484 146076 15540
rect 146132 15484 150000 15540
rect 149200 15456 150000 15484
rect 144274 15260 144284 15316
rect 144340 15260 144956 15316
rect 145012 15260 145022 15316
rect 107762 15036 107772 15092
rect 107828 15036 115836 15092
rect 115892 15036 115902 15092
rect 19612 14868 19622 14924
rect 19678 14868 19726 14924
rect 19782 14868 19830 14924
rect 19886 14868 19896 14924
rect 56432 14868 56442 14924
rect 56498 14868 56546 14924
rect 56602 14868 56650 14924
rect 56706 14868 56716 14924
rect 93252 14868 93262 14924
rect 93318 14868 93366 14924
rect 93422 14868 93470 14924
rect 93526 14868 93536 14924
rect 130072 14868 130082 14924
rect 130138 14868 130186 14924
rect 130242 14868 130290 14924
rect 130346 14868 130356 14924
rect 149200 14644 150000 14672
rect 146066 14588 146076 14644
rect 146132 14588 150000 14644
rect 149200 14560 150000 14588
rect 117394 14364 117404 14420
rect 117460 14364 139468 14420
rect 139524 14364 139534 14420
rect 100482 14252 100492 14308
rect 100548 14252 144396 14308
rect 144452 14252 144956 14308
rect 145012 14252 145022 14308
rect 130498 14140 130508 14196
rect 130564 14140 138572 14196
rect 138628 14140 138638 14196
rect 38022 14084 38032 14140
rect 38088 14084 38136 14140
rect 38192 14084 38240 14140
rect 38296 14084 38306 14140
rect 74842 14084 74852 14140
rect 74908 14084 74956 14140
rect 75012 14084 75060 14140
rect 75116 14084 75126 14140
rect 111662 14084 111672 14140
rect 111728 14084 111776 14140
rect 111832 14084 111880 14140
rect 111936 14084 111946 14140
rect 148482 14084 148492 14140
rect 148548 14084 148596 14140
rect 148652 14084 148700 14140
rect 148756 14084 148766 14140
rect 149200 13748 150000 13776
rect 146066 13692 146076 13748
rect 146132 13692 150000 13748
rect 149200 13664 150000 13692
rect 19612 13300 19622 13356
rect 19678 13300 19726 13356
rect 19782 13300 19830 13356
rect 19886 13300 19896 13356
rect 56432 13300 56442 13356
rect 56498 13300 56546 13356
rect 56602 13300 56650 13356
rect 56706 13300 56716 13356
rect 93252 13300 93262 13356
rect 93318 13300 93366 13356
rect 93422 13300 93470 13356
rect 93526 13300 93536 13356
rect 130072 13300 130082 13356
rect 130138 13300 130186 13356
rect 130242 13300 130290 13356
rect 130346 13300 130356 13356
rect 144386 12908 144396 12964
rect 144452 12908 144956 12964
rect 145012 12908 145022 12964
rect 149200 12852 150000 12880
rect 100034 12796 100044 12852
rect 100100 12796 101164 12852
rect 101220 12796 101230 12852
rect 101490 12796 101500 12852
rect 101556 12796 144284 12852
rect 144340 12796 144350 12852
rect 146066 12796 146076 12852
rect 146132 12796 150000 12852
rect 149200 12768 150000 12796
rect 38022 12516 38032 12572
rect 38088 12516 38136 12572
rect 38192 12516 38240 12572
rect 38296 12516 38306 12572
rect 74842 12516 74852 12572
rect 74908 12516 74956 12572
rect 75012 12516 75060 12572
rect 75116 12516 75126 12572
rect 111662 12516 111672 12572
rect 111728 12516 111776 12572
rect 111832 12516 111880 12572
rect 111936 12516 111946 12572
rect 148482 12516 148492 12572
rect 148548 12516 148596 12572
rect 148652 12516 148700 12572
rect 148756 12516 148766 12572
rect 71362 12348 71372 12404
rect 71428 12348 140028 12404
rect 140084 12348 140094 12404
rect 82786 12236 82796 12292
rect 82852 12236 144620 12292
rect 144676 12236 144686 12292
rect 98466 12124 98476 12180
rect 98532 12124 100156 12180
rect 100212 12124 100222 12180
rect 133522 12012 133532 12068
rect 133588 12012 144284 12068
rect 144340 12012 144956 12068
rect 145012 12012 145022 12068
rect 149200 11956 150000 11984
rect 63858 11900 63868 11956
rect 63924 11900 131964 11956
rect 132020 11900 132030 11956
rect 146066 11900 146076 11956
rect 146132 11900 150000 11956
rect 149200 11872 150000 11900
rect 19612 11732 19622 11788
rect 19678 11732 19726 11788
rect 19782 11732 19830 11788
rect 19886 11732 19896 11788
rect 56432 11732 56442 11788
rect 56498 11732 56546 11788
rect 56602 11732 56650 11788
rect 56706 11732 56716 11788
rect 93252 11732 93262 11788
rect 93318 11732 93366 11788
rect 93422 11732 93470 11788
rect 93526 11732 93536 11788
rect 130072 11732 130082 11788
rect 130138 11732 130186 11788
rect 130242 11732 130290 11788
rect 130346 11732 130356 11788
rect 98018 11116 98028 11172
rect 98084 11116 100492 11172
rect 100548 11116 101164 11172
rect 101220 11116 101230 11172
rect 101490 11116 101500 11172
rect 101556 11116 144284 11172
rect 144340 11116 144350 11172
rect 146066 11116 146076 11172
rect 146132 11116 148932 11172
rect 148876 11060 148932 11116
rect 149200 11060 150000 11088
rect 148876 11004 150000 11060
rect 38022 10948 38032 11004
rect 38088 10948 38136 11004
rect 38192 10948 38240 11004
rect 38296 10948 38306 11004
rect 74842 10948 74852 11004
rect 74908 10948 74956 11004
rect 75012 10948 75060 11004
rect 75116 10948 75126 11004
rect 111662 10948 111672 11004
rect 111728 10948 111776 11004
rect 111832 10948 111880 11004
rect 111936 10948 111946 11004
rect 148482 10948 148492 11004
rect 148548 10948 148596 11004
rect 148652 10948 148700 11004
rect 148756 10948 148766 11004
rect 149200 10976 150000 11004
rect 105858 10780 105868 10836
rect 105924 10780 144396 10836
rect 144452 10780 144956 10836
rect 145012 10780 145022 10836
rect 53890 10668 53900 10724
rect 53956 10668 122108 10724
rect 122164 10668 122174 10724
rect 32386 10556 32396 10612
rect 32452 10556 101948 10612
rect 102004 10556 102014 10612
rect 74722 10444 74732 10500
rect 74788 10444 137564 10500
rect 137620 10444 137630 10500
rect 17042 10332 17052 10388
rect 17108 10332 85596 10388
rect 85652 10332 85662 10388
rect 87154 10332 87164 10388
rect 87220 10332 133980 10388
rect 134036 10332 134046 10388
rect 19612 10164 19622 10220
rect 19678 10164 19726 10220
rect 19782 10164 19830 10220
rect 19886 10164 19896 10220
rect 56432 10164 56442 10220
rect 56498 10164 56546 10220
rect 56602 10164 56650 10220
rect 56706 10164 56716 10220
rect 93252 10164 93262 10220
rect 93318 10164 93366 10220
rect 93422 10164 93470 10220
rect 93526 10164 93536 10220
rect 130072 10164 130082 10220
rect 130138 10164 130186 10220
rect 130242 10164 130290 10220
rect 130346 10164 130356 10220
rect 149200 10164 150000 10192
rect 146290 10108 146300 10164
rect 146356 10108 146860 10164
rect 146916 10108 150000 10164
rect 149200 10080 150000 10108
rect 90738 9884 90748 9940
rect 90804 9884 144956 9940
rect 145012 9884 145022 9940
rect 146290 9660 146300 9716
rect 146356 9660 146972 9716
rect 147028 9660 147038 9716
rect 79426 9548 79436 9604
rect 79492 9548 142716 9604
rect 142772 9548 142782 9604
rect 38022 9380 38032 9436
rect 38088 9380 38136 9436
rect 38192 9380 38240 9436
rect 38296 9380 38306 9436
rect 74842 9380 74852 9436
rect 74908 9380 74956 9436
rect 75012 9380 75060 9436
rect 75116 9380 75126 9436
rect 111662 9380 111672 9436
rect 111728 9380 111776 9436
rect 111832 9380 111880 9436
rect 111936 9380 111946 9436
rect 148482 9380 148492 9436
rect 148548 9380 148596 9436
rect 148652 9380 148700 9436
rect 148756 9380 148766 9436
rect 149200 9268 150000 9296
rect 146962 9212 146972 9268
rect 147028 9212 150000 9268
rect 149200 9184 150000 9212
rect 47170 9100 47180 9156
rect 47236 9100 115276 9156
rect 115332 9100 115342 9156
rect 146290 9100 146300 9156
rect 146356 9100 146860 9156
rect 146916 9100 146926 9156
rect 12114 8988 12124 9044
rect 12180 8988 79772 9044
rect 79828 8988 79838 9044
rect 15026 8876 15036 8932
rect 15092 8876 80668 8932
rect 80724 8876 80734 8932
rect 90290 8876 90300 8932
rect 90356 8876 144956 8932
rect 145012 8876 145022 8932
rect 75618 8764 75628 8820
rect 75684 8764 136220 8820
rect 136276 8764 136286 8820
rect 19612 8596 19622 8652
rect 19678 8596 19726 8652
rect 19782 8596 19830 8652
rect 19886 8596 19896 8652
rect 56432 8596 56442 8652
rect 56498 8596 56546 8652
rect 56602 8596 56650 8652
rect 56706 8596 56716 8652
rect 93252 8596 93262 8652
rect 93318 8596 93366 8652
rect 93422 8596 93470 8652
rect 93526 8596 93536 8652
rect 130072 8596 130082 8652
rect 130138 8596 130186 8652
rect 130242 8596 130290 8652
rect 130346 8596 130356 8652
rect 57026 8428 57036 8484
rect 57092 8428 126924 8484
rect 126980 8428 126990 8484
rect 146850 8428 146860 8484
rect 146916 8428 146926 8484
rect 146860 8372 146916 8428
rect 149200 8372 150000 8400
rect 146860 8316 150000 8372
rect 149200 8288 150000 8316
rect 146290 8092 146300 8148
rect 146356 8092 146972 8148
rect 147028 8092 147038 8148
rect 76178 7980 76188 8036
rect 76244 7980 142716 8036
rect 142772 7980 142782 8036
rect 38022 7812 38032 7868
rect 38088 7812 38136 7868
rect 38192 7812 38240 7868
rect 38296 7812 38306 7868
rect 74842 7812 74852 7868
rect 74908 7812 74956 7868
rect 75012 7812 75060 7868
rect 75116 7812 75126 7868
rect 111662 7812 111672 7868
rect 111728 7812 111776 7868
rect 111832 7812 111880 7868
rect 111936 7812 111946 7868
rect 148482 7812 148492 7868
rect 148548 7812 148596 7868
rect 148652 7812 148700 7868
rect 148756 7812 148766 7868
rect 122658 7756 122668 7812
rect 122724 7756 145068 7812
rect 145124 7756 145134 7812
rect 101490 7644 101500 7700
rect 101556 7644 133532 7700
rect 133588 7644 133598 7700
rect 139906 7644 139916 7700
rect 139972 7644 147084 7700
rect 147140 7644 147150 7700
rect 50978 7532 50988 7588
rect 51044 7532 117964 7588
rect 118020 7532 118030 7588
rect 129826 7532 129836 7588
rect 129892 7532 131292 7588
rect 131348 7532 131740 7588
rect 131796 7532 145180 7588
rect 145236 7532 145246 7588
rect 146178 7532 146188 7588
rect 146244 7532 146860 7588
rect 146916 7532 146926 7588
rect 149200 7476 150000 7504
rect 80546 7420 80556 7476
rect 80612 7420 144956 7476
rect 145012 7420 145022 7476
rect 146962 7420 146972 7476
rect 147028 7420 150000 7476
rect 149200 7392 150000 7420
rect 10770 7308 10780 7364
rect 10836 7308 77980 7364
rect 78036 7308 78046 7364
rect 105522 7308 105532 7364
rect 105588 7308 106652 7364
rect 106708 7308 106718 7364
rect 36306 7196 36316 7252
rect 36372 7196 91532 7252
rect 91588 7196 91598 7252
rect 19612 7028 19622 7084
rect 19678 7028 19726 7084
rect 19782 7028 19830 7084
rect 19886 7028 19896 7084
rect 56432 7028 56442 7084
rect 56498 7028 56546 7084
rect 56602 7028 56650 7084
rect 56706 7028 56716 7084
rect 93252 7028 93262 7084
rect 93318 7028 93366 7084
rect 93422 7028 93470 7084
rect 93526 7028 93536 7084
rect 130072 7028 130082 7084
rect 130138 7028 130186 7084
rect 130242 7028 130290 7084
rect 130346 7028 130356 7084
rect 119298 6972 119308 7028
rect 119364 6972 121772 7028
rect 121828 6972 121838 7028
rect 59826 6860 59836 6916
rect 59892 6860 128828 6916
rect 128884 6860 128894 6916
rect 40338 6748 40348 6804
rect 40404 6748 109116 6804
rect 109172 6748 109182 6804
rect 119186 6748 119196 6804
rect 119252 6748 120204 6804
rect 120260 6748 120270 6804
rect 88386 6636 88396 6692
rect 88452 6636 144732 6692
rect 144788 6636 144798 6692
rect 149200 6580 150000 6608
rect 137554 6524 137564 6580
rect 137620 6524 138124 6580
rect 138180 6524 138190 6580
rect 138898 6524 138908 6580
rect 138964 6524 143164 6580
rect 143220 6524 143230 6580
rect 144274 6524 144284 6580
rect 144340 6524 145180 6580
rect 145236 6524 145246 6580
rect 146290 6524 146300 6580
rect 146356 6524 146972 6580
rect 147028 6524 150000 6580
rect 149200 6496 150000 6524
rect 85652 6412 88900 6468
rect 133634 6412 133644 6468
rect 133700 6412 137004 6468
rect 137060 6412 137788 6468
rect 137844 6412 138684 6468
rect 138740 6412 138750 6468
rect 38022 6244 38032 6300
rect 38088 6244 38136 6300
rect 38192 6244 38240 6300
rect 38296 6244 38306 6300
rect 74842 6244 74852 6300
rect 74908 6244 74956 6300
rect 75012 6244 75060 6300
rect 75116 6244 75126 6300
rect 85652 6244 85708 6412
rect 85362 6188 85372 6244
rect 85428 6188 85708 6244
rect 88844 6244 88900 6412
rect 111662 6244 111672 6300
rect 111728 6244 111776 6300
rect 111832 6244 111880 6300
rect 111936 6244 111946 6300
rect 148482 6244 148492 6300
rect 148548 6244 148596 6300
rect 148652 6244 148700 6300
rect 148756 6244 148766 6300
rect 88844 6188 108388 6244
rect 109106 6188 109116 6244
rect 109172 6188 109900 6244
rect 109956 6188 109966 6244
rect 112028 6188 144956 6244
rect 145012 6188 145022 6244
rect 108332 6132 108388 6188
rect 112028 6132 112084 6188
rect 86930 6076 86940 6132
rect 86996 6076 87836 6132
rect 87892 6076 88396 6132
rect 88452 6076 88462 6132
rect 89180 6076 108276 6132
rect 108332 6076 112084 6132
rect 114212 6076 122668 6132
rect 122724 6076 122734 6132
rect 125972 6076 130340 6132
rect 130498 6076 130508 6132
rect 130564 6076 131068 6132
rect 131124 6076 131134 6132
rect 136210 6076 136220 6132
rect 136276 6076 138236 6132
rect 138292 6076 138302 6132
rect 139682 6076 139692 6132
rect 139748 6076 141148 6132
rect 141204 6076 141214 6132
rect 70578 5964 70588 6020
rect 70644 5964 88956 6020
rect 89012 5964 89022 6020
rect 30034 5852 30044 5908
rect 30100 5852 88956 5908
rect 89012 5852 89022 5908
rect 89180 5796 89236 6076
rect 108220 6020 108276 6076
rect 114212 6020 114268 6076
rect 125972 6020 126028 6076
rect 130284 6020 130340 6076
rect 97346 5964 97356 6020
rect 97412 5964 97916 6020
rect 97972 5964 99036 6020
rect 99092 5964 99102 6020
rect 101938 5964 101948 6020
rect 102004 5964 102732 6020
rect 102788 5964 102798 6020
rect 108220 5964 114268 6020
rect 115266 5964 115276 6020
rect 115332 5964 116060 6020
rect 116116 5964 116126 6020
rect 116498 5964 116508 6020
rect 116564 5964 117740 6020
rect 117796 5964 117806 6020
rect 122098 5964 122108 6020
rect 122164 5964 122892 6020
rect 122948 5964 122958 6020
rect 123116 5964 126028 6020
rect 128818 5964 128828 6020
rect 128884 5964 129500 6020
rect 129556 5964 129566 6020
rect 130284 5964 137788 6020
rect 138674 5964 138684 6020
rect 138740 5964 140364 6020
rect 140420 5964 140430 6020
rect 116508 5908 116564 5964
rect 89394 5852 89404 5908
rect 89460 5852 101388 5908
rect 101444 5852 101454 5908
rect 102162 5852 102172 5908
rect 102228 5852 102620 5908
rect 102676 5852 103740 5908
rect 103796 5852 103806 5908
rect 109778 5852 109788 5908
rect 109844 5852 110460 5908
rect 110516 5852 110526 5908
rect 115378 5852 115388 5908
rect 115444 5852 116564 5908
rect 119074 5852 119084 5908
rect 119140 5852 119756 5908
rect 119812 5852 119822 5908
rect 123116 5796 123172 5964
rect 137732 5908 137788 5964
rect 123890 5852 123900 5908
rect 123956 5852 124572 5908
rect 124628 5852 124638 5908
rect 132626 5852 132636 5908
rect 132692 5852 134428 5908
rect 134484 5852 134494 5908
rect 137732 5852 143500 5908
rect 143556 5852 143566 5908
rect 74498 5740 74508 5796
rect 74564 5740 75740 5796
rect 75796 5740 75806 5796
rect 86034 5740 86044 5796
rect 86100 5740 86940 5796
rect 86996 5740 89236 5796
rect 112018 5740 112028 5796
rect 112084 5740 123172 5796
rect 123330 5740 123340 5796
rect 123396 5740 124348 5796
rect 124404 5740 125468 5796
rect 125524 5740 126588 5796
rect 126644 5740 126654 5796
rect 128930 5740 128940 5796
rect 128996 5740 129948 5796
rect 130004 5740 130956 5796
rect 131012 5740 132076 5796
rect 132132 5740 133756 5796
rect 133812 5740 133822 5796
rect 144050 5740 144060 5796
rect 144116 5740 145964 5796
rect 146020 5740 146860 5796
rect 146916 5740 146926 5796
rect 149200 5684 150000 5712
rect 28578 5628 28588 5684
rect 28644 5628 96460 5684
rect 96516 5628 97468 5684
rect 97524 5628 97534 5684
rect 138898 5628 138908 5684
rect 138964 5628 142940 5684
rect 142996 5628 143006 5684
rect 146290 5628 146300 5684
rect 146356 5628 147308 5684
rect 147364 5628 150000 5684
rect 149200 5600 150000 5628
rect 19612 5460 19622 5516
rect 19678 5460 19726 5516
rect 19782 5460 19830 5516
rect 19886 5460 19896 5516
rect 56432 5460 56442 5516
rect 56498 5460 56546 5516
rect 56602 5460 56650 5516
rect 56706 5460 56716 5516
rect 93252 5460 93262 5516
rect 93318 5460 93366 5516
rect 93422 5460 93470 5516
rect 93526 5460 93536 5516
rect 130072 5460 130082 5516
rect 130138 5460 130186 5516
rect 130242 5460 130290 5516
rect 130346 5460 130356 5516
rect 77186 5404 77196 5460
rect 77252 5404 77644 5460
rect 77700 5404 80556 5460
rect 80612 5404 80622 5460
rect 96012 5404 96460 5460
rect 96516 5404 97020 5460
rect 97076 5404 97086 5460
rect 137330 5404 137340 5460
rect 137396 5404 140924 5460
rect 140980 5404 140990 5460
rect 96012 5348 96068 5404
rect 27122 5292 27132 5348
rect 27188 5292 96068 5348
rect 96226 5292 96236 5348
rect 96292 5292 101164 5348
rect 101220 5292 101230 5348
rect 103730 5292 103740 5348
rect 103796 5292 105868 5348
rect 105924 5292 105934 5348
rect 131730 5292 131740 5348
rect 131796 5292 132972 5348
rect 133028 5292 133038 5348
rect 135426 5292 135436 5348
rect 135492 5292 137004 5348
rect 137060 5292 137070 5348
rect 139234 5292 139244 5348
rect 139300 5292 141820 5348
rect 141876 5292 141886 5348
rect 65650 5180 65660 5236
rect 65716 5180 87164 5236
rect 87220 5180 87230 5236
rect 89394 5180 89404 5236
rect 89460 5180 89852 5236
rect 89908 5180 90188 5236
rect 90244 5180 90748 5236
rect 90804 5180 90814 5236
rect 94098 5180 94108 5236
rect 94164 5180 105644 5236
rect 105700 5180 105710 5236
rect 122322 5180 122332 5236
rect 122388 5180 123452 5236
rect 123508 5180 123518 5236
rect 9986 5068 9996 5124
rect 10052 5068 73836 5124
rect 73892 5068 73902 5124
rect 78530 5068 78540 5124
rect 78596 5068 78876 5124
rect 78932 5068 79436 5124
rect 79492 5068 79502 5124
rect 80994 5068 81004 5124
rect 81060 5068 81452 5124
rect 81508 5068 82236 5124
rect 82292 5068 82796 5124
rect 82852 5068 82862 5124
rect 83346 5068 83356 5124
rect 83412 5068 83804 5124
rect 83860 5068 84588 5124
rect 84644 5068 85372 5124
rect 85428 5068 85438 5124
rect 95442 5068 95452 5124
rect 95508 5068 97132 5124
rect 97188 5068 97198 5124
rect 99250 5068 99260 5124
rect 99316 5068 99484 5124
rect 99540 5068 101052 5124
rect 101108 5068 103852 5124
rect 103908 5068 103918 5124
rect 109554 5068 109564 5124
rect 109620 5068 109788 5124
rect 109844 5068 111468 5124
rect 111524 5068 113148 5124
rect 113204 5068 113214 5124
rect 133522 5068 133532 5124
rect 133588 5068 134652 5124
rect 134708 5068 136556 5124
rect 136612 5068 138460 5124
rect 138516 5068 141148 5124
rect 141204 5068 141214 5124
rect 73378 4956 73388 5012
rect 73444 4956 75404 5012
rect 75460 4956 76188 5012
rect 76244 4956 76254 5012
rect 85474 4956 85484 5012
rect 85540 4956 86044 5012
rect 86100 4956 86110 5012
rect 87714 4956 87724 5012
rect 87780 4956 88172 5012
rect 88228 4956 88238 5012
rect 88946 4956 88956 5012
rect 89012 4956 98588 5012
rect 98644 4956 98924 5012
rect 98980 4956 98990 5012
rect 102452 4956 103964 5012
rect 104020 4956 104412 5012
rect 104468 4956 104478 5012
rect 115714 4956 115724 5012
rect 115780 4956 117180 5012
rect 117236 4956 117246 5012
rect 118290 4956 118300 5012
rect 118356 4956 119868 5012
rect 119924 4956 119934 5012
rect 123106 4956 123116 5012
rect 123172 4956 123788 5012
rect 123844 4956 123854 5012
rect 124898 4956 124908 5012
rect 124964 4956 125132 5012
rect 125188 4956 126812 5012
rect 126868 4956 126878 5012
rect 130834 4956 130844 5012
rect 130900 4956 132972 5012
rect 133028 4956 133308 5012
rect 133364 4956 133374 5012
rect 135874 4956 135884 5012
rect 135940 4956 136444 5012
rect 136500 4956 136510 5012
rect 138338 4956 138348 5012
rect 138404 4956 139804 5012
rect 139860 4956 139870 5012
rect 144610 4956 144620 5012
rect 144676 4956 146860 5012
rect 146916 4956 146926 5012
rect 102452 4900 102508 4956
rect 63746 4844 63756 4900
rect 63812 4844 63980 4900
rect 64036 4844 64316 4900
rect 64372 4844 64382 4900
rect 83906 4844 83916 4900
rect 83972 4844 102508 4900
rect 108322 4844 108332 4900
rect 108388 4844 114268 4900
rect 117058 4844 117068 4900
rect 117124 4844 118972 4900
rect 119028 4844 119038 4900
rect 146290 4844 146300 4900
rect 146356 4844 147420 4900
rect 147476 4844 148932 4900
rect 114212 4788 114268 4844
rect 148876 4788 148932 4844
rect 149200 4788 150000 4816
rect 91522 4732 91532 4788
rect 91588 4732 105644 4788
rect 105700 4732 107100 4788
rect 107156 4732 107166 4788
rect 114212 4732 130620 4788
rect 130676 4732 130686 4788
rect 148876 4732 150000 4788
rect 38022 4676 38032 4732
rect 38088 4676 38136 4732
rect 38192 4676 38240 4732
rect 38296 4676 38306 4732
rect 74842 4676 74852 4732
rect 74908 4676 74956 4732
rect 75012 4676 75060 4732
rect 75116 4676 75126 4732
rect 111662 4676 111672 4732
rect 111728 4676 111776 4732
rect 111832 4676 111880 4732
rect 111936 4676 111946 4732
rect 148482 4676 148492 4732
rect 148548 4676 148596 4732
rect 148652 4676 148700 4732
rect 148756 4676 148766 4732
rect 149200 4704 150000 4732
rect 127586 4620 127596 4676
rect 127652 4620 127932 4676
rect 127988 4620 127998 4676
rect 8754 4508 8764 4564
rect 8820 4508 9772 4564
rect 9828 4508 10780 4564
rect 10836 4508 10846 4564
rect 10994 4508 11004 4564
rect 11060 4508 11340 4564
rect 11396 4508 12124 4564
rect 12180 4508 12190 4564
rect 13010 4508 13020 4564
rect 13076 4508 15036 4564
rect 15092 4508 15102 4564
rect 64082 4508 64092 4564
rect 64148 4508 109228 4564
rect 109284 4508 109294 4564
rect 120194 4508 120204 4564
rect 120260 4508 129276 4564
rect 129332 4508 129342 4564
rect 40786 4396 40796 4452
rect 40852 4396 41692 4452
rect 41748 4396 41758 4452
rect 48850 4396 48860 4452
rect 48916 4396 49644 4452
rect 49700 4396 49710 4452
rect 72594 4396 72604 4452
rect 72660 4396 73500 4452
rect 73556 4396 73566 4452
rect 73826 4396 73836 4452
rect 73892 4396 75628 4452
rect 75684 4396 75694 4452
rect 88274 4396 88284 4452
rect 88340 4396 89292 4452
rect 89348 4396 90300 4452
rect 90356 4396 90366 4452
rect 90514 4396 90524 4452
rect 90580 4396 91084 4452
rect 91140 4396 91150 4452
rect 93986 4396 93996 4452
rect 94052 4396 94220 4452
rect 94276 4396 94556 4452
rect 94612 4396 94622 4452
rect 127810 4396 127820 4452
rect 127876 4396 129164 4452
rect 129220 4396 129230 4452
rect 132850 4396 132860 4452
rect 132916 4396 134428 4452
rect 134484 4396 135772 4452
rect 135828 4396 135838 4452
rect 142146 4396 142156 4452
rect 142212 4396 143836 4452
rect 143892 4396 143902 4452
rect 8306 4284 8316 4340
rect 8372 4284 8876 4340
rect 8932 4284 9996 4340
rect 10052 4284 10062 4340
rect 80098 4284 80108 4340
rect 80164 4284 80556 4340
rect 80612 4284 81452 4340
rect 81508 4284 82124 4340
rect 82180 4284 82190 4340
rect 126802 4284 126812 4340
rect 126868 4284 129276 4340
rect 129332 4284 129342 4340
rect 32946 4172 32956 4228
rect 33012 4172 33740 4228
rect 33796 4172 33806 4228
rect 70690 4172 70700 4228
rect 70756 4172 71820 4228
rect 71876 4172 71886 4228
rect 78978 4172 78988 4228
rect 79044 4172 83020 4228
rect 83076 4172 83086 4228
rect 90850 4172 90860 4228
rect 90916 4172 91756 4228
rect 91812 4172 91822 4228
rect 98242 4172 98252 4228
rect 98308 4172 99036 4228
rect 99092 4172 99102 4228
rect 110898 4172 110908 4228
rect 110964 4172 111804 4228
rect 111860 4172 111870 4228
rect 113810 4172 113820 4228
rect 113876 4172 114380 4228
rect 114436 4172 114446 4228
rect 115378 4172 115388 4228
rect 115444 4172 116060 4228
rect 116116 4172 116126 4228
rect 116722 4172 116732 4228
rect 116788 4172 117516 4228
rect 117572 4172 117582 4228
rect 132290 4172 132300 4228
rect 132356 4172 133420 4228
rect 133476 4172 133486 4228
rect 138114 4172 138124 4228
rect 138180 4172 139020 4228
rect 139076 4172 140028 4228
rect 140084 4172 140094 4228
rect 140802 4172 140812 4228
rect 140868 4172 141820 4228
rect 141876 4172 141886 4228
rect 142034 4172 142044 4228
rect 142100 4172 144956 4228
rect 145012 4172 145022 4228
rect 20066 4060 20076 4116
rect 20132 4060 20524 4116
rect 20580 4060 87388 4116
rect 87444 4060 87454 4116
rect 127586 4060 127596 4116
rect 127652 4060 128492 4116
rect 128548 4060 128558 4116
rect 80770 3948 80780 4004
rect 80836 3948 82684 4004
rect 82740 3948 82750 4004
rect 85652 3948 86380 4004
rect 86436 3948 86446 4004
rect 103282 3948 103292 4004
rect 103348 3948 104300 4004
rect 104356 3948 106316 4004
rect 106372 3948 109564 4004
rect 109620 3948 111020 4004
rect 111076 3948 114268 4004
rect 19612 3892 19622 3948
rect 19678 3892 19726 3948
rect 19782 3892 19830 3948
rect 19886 3892 19896 3948
rect 56432 3892 56442 3948
rect 56498 3892 56546 3948
rect 56602 3892 56650 3948
rect 56706 3892 56716 3948
rect 85652 3892 85708 3948
rect 93252 3892 93262 3948
rect 93318 3892 93366 3948
rect 93422 3892 93470 3948
rect 93526 3892 93536 3948
rect 114212 3892 114268 3948
rect 130072 3892 130082 3948
rect 130138 3892 130186 3948
rect 130242 3892 130290 3948
rect 130346 3892 130356 3948
rect 149200 3892 150000 3920
rect 20626 3836 20636 3892
rect 20692 3836 21420 3892
rect 21476 3836 30492 3892
rect 30548 3836 30558 3892
rect 72706 3836 72716 3892
rect 72772 3836 73388 3892
rect 73444 3836 73454 3892
rect 81788 3836 85708 3892
rect 85810 3836 85820 3892
rect 85876 3836 86716 3892
rect 86772 3836 86782 3892
rect 107426 3836 107436 3892
rect 107492 3836 111188 3892
rect 114212 3836 118076 3892
rect 118132 3836 120204 3892
rect 120260 3836 120270 3892
rect 130946 3836 130956 3892
rect 131012 3836 133644 3892
rect 133700 3836 133710 3892
rect 146290 3836 146300 3892
rect 146356 3836 146860 3892
rect 146916 3836 150000 3892
rect 14914 3724 14924 3780
rect 14980 3724 15148 3780
rect 15204 3724 78988 3780
rect 79044 3724 79054 3780
rect 18274 3612 18284 3668
rect 18340 3612 18732 3668
rect 18788 3612 73108 3668
rect 75730 3612 75740 3668
rect 75796 3612 76972 3668
rect 77028 3612 77038 3668
rect 77410 3612 77420 3668
rect 77476 3612 78764 3668
rect 78820 3612 78830 3668
rect 79090 3612 79100 3668
rect 79156 3612 80892 3668
rect 80948 3612 80958 3668
rect 73052 3556 73108 3612
rect 81788 3556 81844 3836
rect 83244 3724 89068 3780
rect 89124 3724 89134 3780
rect 101378 3724 101388 3780
rect 101444 3724 110908 3780
rect 110964 3724 110974 3780
rect 83244 3668 83300 3724
rect 111132 3668 111188 3836
rect 149200 3808 150000 3836
rect 111346 3724 111356 3780
rect 111412 3724 141148 3780
rect 141204 3724 141484 3780
rect 141540 3724 141550 3780
rect 28690 3500 28700 3556
rect 28756 3500 30268 3556
rect 30324 3500 30334 3556
rect 30482 3500 30492 3556
rect 30548 3500 72436 3556
rect 73052 3500 81844 3556
rect 82236 3612 83300 3668
rect 87490 3612 87500 3668
rect 87556 3612 88732 3668
rect 88788 3612 88798 3668
rect 89170 3612 89180 3668
rect 89236 3612 90524 3668
rect 90580 3612 90590 3668
rect 106418 3612 106428 3668
rect 106484 3612 107660 3668
rect 107716 3612 107726 3668
rect 109330 3612 109340 3668
rect 109396 3612 110908 3668
rect 110964 3612 110974 3668
rect 111132 3612 114268 3668
rect 115826 3612 115836 3668
rect 115892 3612 116732 3668
rect 116788 3612 116798 3668
rect 118738 3612 118748 3668
rect 118804 3612 119644 3668
rect 119700 3612 119710 3668
rect 120642 3612 120652 3668
rect 120708 3612 121548 3668
rect 121604 3612 121614 3668
rect 129266 3612 129276 3668
rect 129332 3612 129836 3668
rect 129892 3612 129902 3668
rect 130498 3612 130508 3668
rect 130564 3612 131180 3668
rect 131236 3612 131246 3668
rect 72380 3444 72436 3500
rect 82236 3444 82292 3612
rect 114212 3556 114268 3612
rect 104290 3500 104300 3556
rect 104356 3500 106204 3556
rect 106260 3500 106764 3556
rect 106820 3500 106830 3556
rect 111010 3500 111020 3556
rect 111076 3500 112588 3556
rect 112644 3500 113484 3556
rect 113540 3500 113550 3556
rect 114212 3500 129332 3556
rect 129490 3500 129500 3556
rect 129556 3500 132188 3556
rect 132244 3500 135324 3556
rect 135380 3500 135390 3556
rect 136210 3500 136220 3556
rect 136276 3500 137004 3556
rect 137060 3500 137788 3556
rect 129276 3444 129332 3500
rect 137732 3444 137788 3500
rect 5170 3388 5180 3444
rect 5236 3388 5852 3444
rect 5908 3388 5918 3444
rect 23650 3388 23660 3444
rect 23716 3388 25228 3444
rect 25284 3388 25294 3444
rect 27122 3388 27132 3444
rect 27188 3388 29148 3444
rect 29204 3388 29214 3444
rect 31378 3388 31388 3444
rect 31444 3388 32060 3444
rect 32116 3388 33068 3444
rect 33124 3388 33134 3444
rect 35410 3388 35420 3444
rect 35476 3388 36988 3444
rect 37044 3388 37054 3444
rect 38882 3388 38892 3444
rect 38948 3388 40908 3444
rect 40964 3388 40974 3444
rect 43810 3388 43820 3444
rect 43876 3388 45388 3444
rect 45444 3388 45454 3444
rect 47170 3388 47180 3444
rect 47236 3388 48748 3444
rect 48804 3388 48814 3444
rect 50642 3388 50652 3444
rect 50708 3388 52668 3444
rect 52724 3388 52734 3444
rect 58930 3388 58940 3444
rect 58996 3388 60508 3444
rect 60564 3388 60574 3444
rect 62402 3388 62412 3444
rect 62468 3388 64428 3444
rect 64484 3388 64494 3444
rect 67330 3388 67340 3444
rect 67396 3388 68908 3444
rect 68964 3388 68974 3444
rect 72380 3388 82292 3444
rect 82450 3388 82460 3444
rect 82516 3388 83356 3444
rect 83412 3388 83422 3444
rect 95218 3388 95228 3444
rect 95284 3388 95900 3444
rect 95956 3388 96236 3444
rect 96292 3388 96302 3444
rect 97570 3388 97580 3444
rect 97636 3388 98028 3444
rect 98084 3388 98094 3444
rect 99250 3388 99260 3444
rect 99316 3388 100828 3444
rect 100884 3388 100894 3444
rect 103058 3388 103068 3444
rect 103124 3388 104748 3444
rect 104804 3388 104814 3444
rect 105970 3388 105980 3444
rect 106036 3388 107884 3444
rect 107940 3388 108668 3444
rect 108724 3388 108734 3444
rect 112690 3388 112700 3444
rect 112756 3388 113260 3444
rect 113316 3388 113932 3444
rect 113988 3388 113998 3444
rect 114818 3388 114828 3444
rect 114884 3388 115612 3444
rect 115668 3388 115678 3444
rect 117730 3388 117740 3444
rect 117796 3388 118524 3444
rect 118580 3388 119196 3444
rect 119252 3388 119262 3444
rect 119410 3388 119420 3444
rect 119476 3388 120652 3444
rect 120708 3388 120718 3444
rect 121090 3388 121100 3444
rect 121156 3388 121436 3444
rect 121492 3388 121996 3444
rect 122052 3388 122062 3444
rect 122770 3388 122780 3444
rect 122836 3388 124348 3444
rect 124404 3388 124414 3444
rect 126130 3388 126140 3444
rect 126196 3388 127372 3444
rect 127428 3388 127438 3444
rect 129276 3388 130956 3444
rect 131012 3388 131022 3444
rect 131170 3388 131180 3444
rect 131236 3388 132412 3444
rect 132468 3388 134204 3444
rect 134260 3388 134270 3444
rect 134530 3388 134540 3444
rect 134596 3388 136108 3444
rect 136164 3388 136174 3444
rect 137732 3388 138012 3444
rect 138068 3388 138078 3444
rect 139570 3388 139580 3444
rect 139636 3388 140140 3444
rect 140196 3388 140924 3444
rect 140980 3388 140990 3444
rect 141250 3388 141260 3444
rect 141316 3388 141820 3444
rect 141876 3388 142716 3444
rect 142772 3388 142782 3444
rect 142930 3388 142940 3444
rect 142996 3388 144172 3444
rect 144228 3388 145068 3444
rect 145124 3388 145134 3444
rect 6962 3276 6972 3332
rect 7028 3276 73164 3332
rect 73220 3276 73230 3332
rect 85586 3276 85596 3332
rect 85652 3276 86156 3332
rect 86212 3276 86222 3332
rect 138226 3276 138236 3332
rect 138292 3276 147868 3332
rect 147924 3276 147934 3332
rect 38022 3108 38032 3164
rect 38088 3108 38136 3164
rect 38192 3108 38240 3164
rect 38296 3108 38306 3164
rect 74842 3108 74852 3164
rect 74908 3108 74956 3164
rect 75012 3108 75060 3164
rect 75116 3108 75126 3164
rect 111662 3108 111672 3164
rect 111728 3108 111776 3164
rect 111832 3108 111880 3164
rect 111936 3108 111946 3164
rect 148482 3108 148492 3164
rect 148548 3108 148596 3164
rect 148652 3108 148700 3164
rect 148756 3108 148766 3164
rect 149200 2996 150000 3024
rect 55458 2940 55468 2996
rect 55524 2940 124908 2996
rect 124964 2940 124974 2996
rect 145170 2940 145180 2996
rect 145236 2940 150000 2996
rect 149200 2912 150000 2940
rect 43026 2828 43036 2884
rect 43092 2828 111132 2884
rect 111188 2828 112252 2884
rect 112308 2828 112318 2884
rect 48066 2716 48076 2772
rect 48132 2716 115724 2772
rect 115780 2716 115790 2772
rect 38658 2604 38668 2660
rect 38724 2604 64092 2660
rect 64148 2604 64158 2660
rect 82114 2604 82124 2660
rect 82180 2604 142044 2660
rect 142100 2604 142110 2660
rect 62178 2492 62188 2548
rect 62244 2492 108332 2548
rect 108388 2492 108398 2548
rect 110674 2492 110684 2548
rect 110740 2492 143948 2548
rect 144004 2492 144014 2548
rect 23762 2380 23772 2436
rect 23828 2380 106092 2436
rect 106148 2380 106158 2436
rect 31938 2268 31948 2324
rect 32004 2268 101836 2324
rect 101892 2268 101902 2324
rect 149200 2100 150000 2128
rect 146066 2044 146076 2100
rect 146132 2044 150000 2100
rect 149200 2016 150000 2044
rect 24546 1596 24556 1652
rect 24612 1596 94668 1652
rect 94724 1596 94734 1652
rect 45154 1484 45164 1540
rect 45220 1484 115052 1540
rect 115108 1484 115118 1540
rect 68674 1372 68684 1428
rect 68740 1372 138348 1428
rect 138404 1372 138414 1428
rect 52098 1260 52108 1316
rect 52164 1260 121324 1316
rect 121380 1260 121390 1316
rect 149200 1204 150000 1232
rect 59042 1148 59052 1204
rect 59108 1148 128828 1204
rect 128884 1148 128894 1204
rect 145954 1148 145964 1204
rect 146020 1148 150000 1204
rect 149200 1120 150000 1148
rect 43698 1036 43708 1092
rect 43764 1036 113036 1092
rect 113092 1036 113102 1092
rect 67218 924 67228 980
rect 67284 924 136444 980
rect 136500 924 136510 980
rect 35634 812 35644 868
rect 35700 812 83916 868
rect 83972 812 83982 868
<< via3 >>
rect 19622 36820 19678 36876
rect 19726 36820 19782 36876
rect 19830 36820 19886 36876
rect 56442 36820 56498 36876
rect 56546 36820 56602 36876
rect 56650 36820 56706 36876
rect 93262 36820 93318 36876
rect 93366 36820 93422 36876
rect 93470 36820 93526 36876
rect 130082 36820 130138 36876
rect 130186 36820 130242 36876
rect 130290 36820 130346 36876
rect 38032 36036 38088 36092
rect 38136 36036 38192 36092
rect 38240 36036 38296 36092
rect 74852 36036 74908 36092
rect 74956 36036 75012 36092
rect 75060 36036 75116 36092
rect 111672 36036 111728 36092
rect 111776 36036 111832 36092
rect 111880 36036 111936 36092
rect 148492 36036 148548 36092
rect 148596 36036 148652 36092
rect 148700 36036 148756 36092
rect 19622 35252 19678 35308
rect 19726 35252 19782 35308
rect 19830 35252 19886 35308
rect 56442 35252 56498 35308
rect 56546 35252 56602 35308
rect 56650 35252 56706 35308
rect 93262 35252 93318 35308
rect 93366 35252 93422 35308
rect 93470 35252 93526 35308
rect 130082 35252 130138 35308
rect 130186 35252 130242 35308
rect 130290 35252 130346 35308
rect 38032 34468 38088 34524
rect 38136 34468 38192 34524
rect 38240 34468 38296 34524
rect 74852 34468 74908 34524
rect 74956 34468 75012 34524
rect 75060 34468 75116 34524
rect 111672 34468 111728 34524
rect 111776 34468 111832 34524
rect 111880 34468 111936 34524
rect 148492 34468 148548 34524
rect 148596 34468 148652 34524
rect 148700 34468 148756 34524
rect 19622 33684 19678 33740
rect 19726 33684 19782 33740
rect 19830 33684 19886 33740
rect 56442 33684 56498 33740
rect 56546 33684 56602 33740
rect 56650 33684 56706 33740
rect 93262 33684 93318 33740
rect 93366 33684 93422 33740
rect 93470 33684 93526 33740
rect 130082 33684 130138 33740
rect 130186 33684 130242 33740
rect 130290 33684 130346 33740
rect 38032 32900 38088 32956
rect 38136 32900 38192 32956
rect 38240 32900 38296 32956
rect 74852 32900 74908 32956
rect 74956 32900 75012 32956
rect 75060 32900 75116 32956
rect 111672 32900 111728 32956
rect 111776 32900 111832 32956
rect 111880 32900 111936 32956
rect 148492 32900 148548 32956
rect 148596 32900 148652 32956
rect 148700 32900 148756 32956
rect 19622 32116 19678 32172
rect 19726 32116 19782 32172
rect 19830 32116 19886 32172
rect 56442 32116 56498 32172
rect 56546 32116 56602 32172
rect 56650 32116 56706 32172
rect 93262 32116 93318 32172
rect 93366 32116 93422 32172
rect 93470 32116 93526 32172
rect 130082 32116 130138 32172
rect 130186 32116 130242 32172
rect 130290 32116 130346 32172
rect 38032 31332 38088 31388
rect 38136 31332 38192 31388
rect 38240 31332 38296 31388
rect 74852 31332 74908 31388
rect 74956 31332 75012 31388
rect 75060 31332 75116 31388
rect 111672 31332 111728 31388
rect 111776 31332 111832 31388
rect 111880 31332 111936 31388
rect 148492 31332 148548 31388
rect 148596 31332 148652 31388
rect 148700 31332 148756 31388
rect 19622 30548 19678 30604
rect 19726 30548 19782 30604
rect 19830 30548 19886 30604
rect 56442 30548 56498 30604
rect 56546 30548 56602 30604
rect 56650 30548 56706 30604
rect 93262 30548 93318 30604
rect 93366 30548 93422 30604
rect 93470 30548 93526 30604
rect 130082 30548 130138 30604
rect 130186 30548 130242 30604
rect 130290 30548 130346 30604
rect 38032 29764 38088 29820
rect 38136 29764 38192 29820
rect 38240 29764 38296 29820
rect 74852 29764 74908 29820
rect 74956 29764 75012 29820
rect 75060 29764 75116 29820
rect 111672 29764 111728 29820
rect 111776 29764 111832 29820
rect 111880 29764 111936 29820
rect 148492 29764 148548 29820
rect 148596 29764 148652 29820
rect 148700 29764 148756 29820
rect 19622 28980 19678 29036
rect 19726 28980 19782 29036
rect 19830 28980 19886 29036
rect 56442 28980 56498 29036
rect 56546 28980 56602 29036
rect 56650 28980 56706 29036
rect 93262 28980 93318 29036
rect 93366 28980 93422 29036
rect 93470 28980 93526 29036
rect 130082 28980 130138 29036
rect 130186 28980 130242 29036
rect 130290 28980 130346 29036
rect 38032 28196 38088 28252
rect 38136 28196 38192 28252
rect 38240 28196 38296 28252
rect 74852 28196 74908 28252
rect 74956 28196 75012 28252
rect 75060 28196 75116 28252
rect 111672 28196 111728 28252
rect 111776 28196 111832 28252
rect 111880 28196 111936 28252
rect 148492 28196 148548 28252
rect 148596 28196 148652 28252
rect 148700 28196 148756 28252
rect 19622 27412 19678 27468
rect 19726 27412 19782 27468
rect 19830 27412 19886 27468
rect 56442 27412 56498 27468
rect 56546 27412 56602 27468
rect 56650 27412 56706 27468
rect 93262 27412 93318 27468
rect 93366 27412 93422 27468
rect 93470 27412 93526 27468
rect 130082 27412 130138 27468
rect 130186 27412 130242 27468
rect 130290 27412 130346 27468
rect 38032 26628 38088 26684
rect 38136 26628 38192 26684
rect 38240 26628 38296 26684
rect 74852 26628 74908 26684
rect 74956 26628 75012 26684
rect 75060 26628 75116 26684
rect 111672 26628 111728 26684
rect 111776 26628 111832 26684
rect 111880 26628 111936 26684
rect 148492 26628 148548 26684
rect 148596 26628 148652 26684
rect 148700 26628 148756 26684
rect 19622 25844 19678 25900
rect 19726 25844 19782 25900
rect 19830 25844 19886 25900
rect 56442 25844 56498 25900
rect 56546 25844 56602 25900
rect 56650 25844 56706 25900
rect 93262 25844 93318 25900
rect 93366 25844 93422 25900
rect 93470 25844 93526 25900
rect 130082 25844 130138 25900
rect 130186 25844 130242 25900
rect 130290 25844 130346 25900
rect 38032 25060 38088 25116
rect 38136 25060 38192 25116
rect 38240 25060 38296 25116
rect 74852 25060 74908 25116
rect 74956 25060 75012 25116
rect 75060 25060 75116 25116
rect 111672 25060 111728 25116
rect 111776 25060 111832 25116
rect 111880 25060 111936 25116
rect 148492 25060 148548 25116
rect 148596 25060 148652 25116
rect 148700 25060 148756 25116
rect 19622 24276 19678 24332
rect 19726 24276 19782 24332
rect 19830 24276 19886 24332
rect 56442 24276 56498 24332
rect 56546 24276 56602 24332
rect 56650 24276 56706 24332
rect 93262 24276 93318 24332
rect 93366 24276 93422 24332
rect 93470 24276 93526 24332
rect 130082 24276 130138 24332
rect 130186 24276 130242 24332
rect 130290 24276 130346 24332
rect 38032 23492 38088 23548
rect 38136 23492 38192 23548
rect 38240 23492 38296 23548
rect 74852 23492 74908 23548
rect 74956 23492 75012 23548
rect 75060 23492 75116 23548
rect 111672 23492 111728 23548
rect 111776 23492 111832 23548
rect 111880 23492 111936 23548
rect 148492 23492 148548 23548
rect 148596 23492 148652 23548
rect 148700 23492 148756 23548
rect 19622 22708 19678 22764
rect 19726 22708 19782 22764
rect 19830 22708 19886 22764
rect 56442 22708 56498 22764
rect 56546 22708 56602 22764
rect 56650 22708 56706 22764
rect 93262 22708 93318 22764
rect 93366 22708 93422 22764
rect 93470 22708 93526 22764
rect 130082 22708 130138 22764
rect 130186 22708 130242 22764
rect 130290 22708 130346 22764
rect 38032 21924 38088 21980
rect 38136 21924 38192 21980
rect 38240 21924 38296 21980
rect 74852 21924 74908 21980
rect 74956 21924 75012 21980
rect 75060 21924 75116 21980
rect 111672 21924 111728 21980
rect 111776 21924 111832 21980
rect 111880 21924 111936 21980
rect 148492 21924 148548 21980
rect 148596 21924 148652 21980
rect 148700 21924 148756 21980
rect 19622 21140 19678 21196
rect 19726 21140 19782 21196
rect 19830 21140 19886 21196
rect 56442 21140 56498 21196
rect 56546 21140 56602 21196
rect 56650 21140 56706 21196
rect 93262 21140 93318 21196
rect 93366 21140 93422 21196
rect 93470 21140 93526 21196
rect 130082 21140 130138 21196
rect 130186 21140 130242 21196
rect 130290 21140 130346 21196
rect 38032 20356 38088 20412
rect 38136 20356 38192 20412
rect 38240 20356 38296 20412
rect 74852 20356 74908 20412
rect 74956 20356 75012 20412
rect 75060 20356 75116 20412
rect 111672 20356 111728 20412
rect 111776 20356 111832 20412
rect 111880 20356 111936 20412
rect 148492 20356 148548 20412
rect 148596 20356 148652 20412
rect 148700 20356 148756 20412
rect 19622 19572 19678 19628
rect 19726 19572 19782 19628
rect 19830 19572 19886 19628
rect 56442 19572 56498 19628
rect 56546 19572 56602 19628
rect 56650 19572 56706 19628
rect 93262 19572 93318 19628
rect 93366 19572 93422 19628
rect 93470 19572 93526 19628
rect 130082 19572 130138 19628
rect 130186 19572 130242 19628
rect 130290 19572 130346 19628
rect 38032 18788 38088 18844
rect 38136 18788 38192 18844
rect 38240 18788 38296 18844
rect 74852 18788 74908 18844
rect 74956 18788 75012 18844
rect 75060 18788 75116 18844
rect 111672 18788 111728 18844
rect 111776 18788 111832 18844
rect 111880 18788 111936 18844
rect 148492 18788 148548 18844
rect 148596 18788 148652 18844
rect 148700 18788 148756 18844
rect 19622 18004 19678 18060
rect 19726 18004 19782 18060
rect 19830 18004 19886 18060
rect 56442 18004 56498 18060
rect 56546 18004 56602 18060
rect 56650 18004 56706 18060
rect 93262 18004 93318 18060
rect 93366 18004 93422 18060
rect 93470 18004 93526 18060
rect 130082 18004 130138 18060
rect 130186 18004 130242 18060
rect 130290 18004 130346 18060
rect 38032 17220 38088 17276
rect 38136 17220 38192 17276
rect 38240 17220 38296 17276
rect 74852 17220 74908 17276
rect 74956 17220 75012 17276
rect 75060 17220 75116 17276
rect 111672 17220 111728 17276
rect 111776 17220 111832 17276
rect 111880 17220 111936 17276
rect 148492 17220 148548 17276
rect 148596 17220 148652 17276
rect 148700 17220 148756 17276
rect 19622 16436 19678 16492
rect 19726 16436 19782 16492
rect 19830 16436 19886 16492
rect 56442 16436 56498 16492
rect 56546 16436 56602 16492
rect 56650 16436 56706 16492
rect 93262 16436 93318 16492
rect 93366 16436 93422 16492
rect 93470 16436 93526 16492
rect 130082 16436 130138 16492
rect 130186 16436 130242 16492
rect 130290 16436 130346 16492
rect 38032 15652 38088 15708
rect 38136 15652 38192 15708
rect 38240 15652 38296 15708
rect 74852 15652 74908 15708
rect 74956 15652 75012 15708
rect 75060 15652 75116 15708
rect 111672 15652 111728 15708
rect 111776 15652 111832 15708
rect 111880 15652 111936 15708
rect 148492 15652 148548 15708
rect 148596 15652 148652 15708
rect 148700 15652 148756 15708
rect 19622 14868 19678 14924
rect 19726 14868 19782 14924
rect 19830 14868 19886 14924
rect 56442 14868 56498 14924
rect 56546 14868 56602 14924
rect 56650 14868 56706 14924
rect 93262 14868 93318 14924
rect 93366 14868 93422 14924
rect 93470 14868 93526 14924
rect 130082 14868 130138 14924
rect 130186 14868 130242 14924
rect 130290 14868 130346 14924
rect 38032 14084 38088 14140
rect 38136 14084 38192 14140
rect 38240 14084 38296 14140
rect 74852 14084 74908 14140
rect 74956 14084 75012 14140
rect 75060 14084 75116 14140
rect 111672 14084 111728 14140
rect 111776 14084 111832 14140
rect 111880 14084 111936 14140
rect 148492 14084 148548 14140
rect 148596 14084 148652 14140
rect 148700 14084 148756 14140
rect 19622 13300 19678 13356
rect 19726 13300 19782 13356
rect 19830 13300 19886 13356
rect 56442 13300 56498 13356
rect 56546 13300 56602 13356
rect 56650 13300 56706 13356
rect 93262 13300 93318 13356
rect 93366 13300 93422 13356
rect 93470 13300 93526 13356
rect 130082 13300 130138 13356
rect 130186 13300 130242 13356
rect 130290 13300 130346 13356
rect 38032 12516 38088 12572
rect 38136 12516 38192 12572
rect 38240 12516 38296 12572
rect 74852 12516 74908 12572
rect 74956 12516 75012 12572
rect 75060 12516 75116 12572
rect 111672 12516 111728 12572
rect 111776 12516 111832 12572
rect 111880 12516 111936 12572
rect 148492 12516 148548 12572
rect 148596 12516 148652 12572
rect 148700 12516 148756 12572
rect 19622 11732 19678 11788
rect 19726 11732 19782 11788
rect 19830 11732 19886 11788
rect 56442 11732 56498 11788
rect 56546 11732 56602 11788
rect 56650 11732 56706 11788
rect 93262 11732 93318 11788
rect 93366 11732 93422 11788
rect 93470 11732 93526 11788
rect 130082 11732 130138 11788
rect 130186 11732 130242 11788
rect 130290 11732 130346 11788
rect 38032 10948 38088 11004
rect 38136 10948 38192 11004
rect 38240 10948 38296 11004
rect 74852 10948 74908 11004
rect 74956 10948 75012 11004
rect 75060 10948 75116 11004
rect 111672 10948 111728 11004
rect 111776 10948 111832 11004
rect 111880 10948 111936 11004
rect 148492 10948 148548 11004
rect 148596 10948 148652 11004
rect 148700 10948 148756 11004
rect 19622 10164 19678 10220
rect 19726 10164 19782 10220
rect 19830 10164 19886 10220
rect 56442 10164 56498 10220
rect 56546 10164 56602 10220
rect 56650 10164 56706 10220
rect 93262 10164 93318 10220
rect 93366 10164 93422 10220
rect 93470 10164 93526 10220
rect 130082 10164 130138 10220
rect 130186 10164 130242 10220
rect 130290 10164 130346 10220
rect 38032 9380 38088 9436
rect 38136 9380 38192 9436
rect 38240 9380 38296 9436
rect 74852 9380 74908 9436
rect 74956 9380 75012 9436
rect 75060 9380 75116 9436
rect 111672 9380 111728 9436
rect 111776 9380 111832 9436
rect 111880 9380 111936 9436
rect 148492 9380 148548 9436
rect 148596 9380 148652 9436
rect 148700 9380 148756 9436
rect 19622 8596 19678 8652
rect 19726 8596 19782 8652
rect 19830 8596 19886 8652
rect 56442 8596 56498 8652
rect 56546 8596 56602 8652
rect 56650 8596 56706 8652
rect 93262 8596 93318 8652
rect 93366 8596 93422 8652
rect 93470 8596 93526 8652
rect 130082 8596 130138 8652
rect 130186 8596 130242 8652
rect 130290 8596 130346 8652
rect 38032 7812 38088 7868
rect 38136 7812 38192 7868
rect 38240 7812 38296 7868
rect 74852 7812 74908 7868
rect 74956 7812 75012 7868
rect 75060 7812 75116 7868
rect 111672 7812 111728 7868
rect 111776 7812 111832 7868
rect 111880 7812 111936 7868
rect 148492 7812 148548 7868
rect 148596 7812 148652 7868
rect 148700 7812 148756 7868
rect 19622 7028 19678 7084
rect 19726 7028 19782 7084
rect 19830 7028 19886 7084
rect 56442 7028 56498 7084
rect 56546 7028 56602 7084
rect 56650 7028 56706 7084
rect 93262 7028 93318 7084
rect 93366 7028 93422 7084
rect 93470 7028 93526 7084
rect 130082 7028 130138 7084
rect 130186 7028 130242 7084
rect 130290 7028 130346 7084
rect 38032 6244 38088 6300
rect 38136 6244 38192 6300
rect 38240 6244 38296 6300
rect 74852 6244 74908 6300
rect 74956 6244 75012 6300
rect 75060 6244 75116 6300
rect 111672 6244 111728 6300
rect 111776 6244 111832 6300
rect 111880 6244 111936 6300
rect 148492 6244 148548 6300
rect 148596 6244 148652 6300
rect 148700 6244 148756 6300
rect 88956 5964 89012 6020
rect 89404 5852 89460 5908
rect 19622 5460 19678 5516
rect 19726 5460 19782 5516
rect 19830 5460 19886 5516
rect 56442 5460 56498 5516
rect 56546 5460 56602 5516
rect 56650 5460 56706 5516
rect 93262 5460 93318 5516
rect 93366 5460 93422 5516
rect 93470 5460 93526 5516
rect 130082 5460 130138 5516
rect 130186 5460 130242 5516
rect 130290 5460 130346 5516
rect 38032 4676 38088 4732
rect 38136 4676 38192 4732
rect 38240 4676 38296 4732
rect 74852 4676 74908 4732
rect 74956 4676 75012 4732
rect 75060 4676 75116 4732
rect 111672 4676 111728 4732
rect 111776 4676 111832 4732
rect 111880 4676 111936 4732
rect 148492 4676 148548 4732
rect 148596 4676 148652 4732
rect 148700 4676 148756 4732
rect 19622 3892 19678 3948
rect 19726 3892 19782 3948
rect 19830 3892 19886 3948
rect 56442 3892 56498 3948
rect 56546 3892 56602 3948
rect 56650 3892 56706 3948
rect 93262 3892 93318 3948
rect 93366 3892 93422 3948
rect 93470 3892 93526 3948
rect 130082 3892 130138 3948
rect 130186 3892 130242 3948
rect 130290 3892 130346 3948
rect 30492 3836 30548 3892
rect 130956 3836 131012 3892
rect 110908 3724 110964 3780
rect 111356 3724 111412 3780
rect 30492 3500 30548 3556
rect 130956 3388 131012 3444
rect 38032 3108 38088 3164
rect 38136 3108 38192 3164
rect 38240 3108 38296 3164
rect 74852 3108 74908 3164
rect 74956 3108 75012 3164
rect 75060 3108 75116 3164
rect 111672 3108 111728 3164
rect 111776 3108 111832 3164
rect 111880 3108 111936 3164
rect 148492 3108 148548 3164
rect 148596 3108 148652 3164
rect 148700 3108 148756 3164
<< metal4 >>
rect 19594 36876 19914 36908
rect 19594 36820 19622 36876
rect 19678 36820 19726 36876
rect 19782 36820 19830 36876
rect 19886 36820 19914 36876
rect 19594 35308 19914 36820
rect 19594 35252 19622 35308
rect 19678 35252 19726 35308
rect 19782 35252 19830 35308
rect 19886 35252 19914 35308
rect 19594 33740 19914 35252
rect 19594 33684 19622 33740
rect 19678 33684 19726 33740
rect 19782 33684 19830 33740
rect 19886 33684 19914 33740
rect 19594 32172 19914 33684
rect 19594 32116 19622 32172
rect 19678 32116 19726 32172
rect 19782 32116 19830 32172
rect 19886 32116 19914 32172
rect 19594 30604 19914 32116
rect 19594 30548 19622 30604
rect 19678 30548 19726 30604
rect 19782 30548 19830 30604
rect 19886 30548 19914 30604
rect 19594 29036 19914 30548
rect 19594 28980 19622 29036
rect 19678 28980 19726 29036
rect 19782 28980 19830 29036
rect 19886 28980 19914 29036
rect 19594 27468 19914 28980
rect 19594 27412 19622 27468
rect 19678 27412 19726 27468
rect 19782 27412 19830 27468
rect 19886 27412 19914 27468
rect 19594 25900 19914 27412
rect 19594 25844 19622 25900
rect 19678 25844 19726 25900
rect 19782 25844 19830 25900
rect 19886 25844 19914 25900
rect 19594 24332 19914 25844
rect 19594 24276 19622 24332
rect 19678 24276 19726 24332
rect 19782 24276 19830 24332
rect 19886 24276 19914 24332
rect 19594 22764 19914 24276
rect 19594 22708 19622 22764
rect 19678 22708 19726 22764
rect 19782 22708 19830 22764
rect 19886 22708 19914 22764
rect 19594 21196 19914 22708
rect 19594 21140 19622 21196
rect 19678 21140 19726 21196
rect 19782 21140 19830 21196
rect 19886 21140 19914 21196
rect 19594 19628 19914 21140
rect 19594 19572 19622 19628
rect 19678 19572 19726 19628
rect 19782 19572 19830 19628
rect 19886 19572 19914 19628
rect 19594 18060 19914 19572
rect 19594 18004 19622 18060
rect 19678 18004 19726 18060
rect 19782 18004 19830 18060
rect 19886 18004 19914 18060
rect 19594 16492 19914 18004
rect 19594 16436 19622 16492
rect 19678 16436 19726 16492
rect 19782 16436 19830 16492
rect 19886 16436 19914 16492
rect 19594 14924 19914 16436
rect 19594 14868 19622 14924
rect 19678 14868 19726 14924
rect 19782 14868 19830 14924
rect 19886 14868 19914 14924
rect 19594 13356 19914 14868
rect 19594 13300 19622 13356
rect 19678 13300 19726 13356
rect 19782 13300 19830 13356
rect 19886 13300 19914 13356
rect 19594 11788 19914 13300
rect 19594 11732 19622 11788
rect 19678 11732 19726 11788
rect 19782 11732 19830 11788
rect 19886 11732 19914 11788
rect 19594 10220 19914 11732
rect 19594 10164 19622 10220
rect 19678 10164 19726 10220
rect 19782 10164 19830 10220
rect 19886 10164 19914 10220
rect 19594 8652 19914 10164
rect 19594 8596 19622 8652
rect 19678 8596 19726 8652
rect 19782 8596 19830 8652
rect 19886 8596 19914 8652
rect 19594 7084 19914 8596
rect 19594 7028 19622 7084
rect 19678 7028 19726 7084
rect 19782 7028 19830 7084
rect 19886 7028 19914 7084
rect 19594 5516 19914 7028
rect 19594 5460 19622 5516
rect 19678 5460 19726 5516
rect 19782 5460 19830 5516
rect 19886 5460 19914 5516
rect 19594 3948 19914 5460
rect 19594 3892 19622 3948
rect 19678 3892 19726 3948
rect 19782 3892 19830 3948
rect 19886 3892 19914 3948
rect 38004 36092 38324 36908
rect 38004 36036 38032 36092
rect 38088 36036 38136 36092
rect 38192 36036 38240 36092
rect 38296 36036 38324 36092
rect 38004 34524 38324 36036
rect 38004 34468 38032 34524
rect 38088 34468 38136 34524
rect 38192 34468 38240 34524
rect 38296 34468 38324 34524
rect 38004 32956 38324 34468
rect 38004 32900 38032 32956
rect 38088 32900 38136 32956
rect 38192 32900 38240 32956
rect 38296 32900 38324 32956
rect 38004 31388 38324 32900
rect 38004 31332 38032 31388
rect 38088 31332 38136 31388
rect 38192 31332 38240 31388
rect 38296 31332 38324 31388
rect 38004 29820 38324 31332
rect 38004 29764 38032 29820
rect 38088 29764 38136 29820
rect 38192 29764 38240 29820
rect 38296 29764 38324 29820
rect 38004 28252 38324 29764
rect 38004 28196 38032 28252
rect 38088 28196 38136 28252
rect 38192 28196 38240 28252
rect 38296 28196 38324 28252
rect 38004 26684 38324 28196
rect 38004 26628 38032 26684
rect 38088 26628 38136 26684
rect 38192 26628 38240 26684
rect 38296 26628 38324 26684
rect 38004 25116 38324 26628
rect 38004 25060 38032 25116
rect 38088 25060 38136 25116
rect 38192 25060 38240 25116
rect 38296 25060 38324 25116
rect 38004 23548 38324 25060
rect 38004 23492 38032 23548
rect 38088 23492 38136 23548
rect 38192 23492 38240 23548
rect 38296 23492 38324 23548
rect 38004 21980 38324 23492
rect 38004 21924 38032 21980
rect 38088 21924 38136 21980
rect 38192 21924 38240 21980
rect 38296 21924 38324 21980
rect 38004 20412 38324 21924
rect 38004 20356 38032 20412
rect 38088 20356 38136 20412
rect 38192 20356 38240 20412
rect 38296 20356 38324 20412
rect 38004 18844 38324 20356
rect 38004 18788 38032 18844
rect 38088 18788 38136 18844
rect 38192 18788 38240 18844
rect 38296 18788 38324 18844
rect 38004 17276 38324 18788
rect 38004 17220 38032 17276
rect 38088 17220 38136 17276
rect 38192 17220 38240 17276
rect 38296 17220 38324 17276
rect 38004 15708 38324 17220
rect 38004 15652 38032 15708
rect 38088 15652 38136 15708
rect 38192 15652 38240 15708
rect 38296 15652 38324 15708
rect 38004 14140 38324 15652
rect 38004 14084 38032 14140
rect 38088 14084 38136 14140
rect 38192 14084 38240 14140
rect 38296 14084 38324 14140
rect 38004 12572 38324 14084
rect 38004 12516 38032 12572
rect 38088 12516 38136 12572
rect 38192 12516 38240 12572
rect 38296 12516 38324 12572
rect 38004 11004 38324 12516
rect 38004 10948 38032 11004
rect 38088 10948 38136 11004
rect 38192 10948 38240 11004
rect 38296 10948 38324 11004
rect 38004 9436 38324 10948
rect 38004 9380 38032 9436
rect 38088 9380 38136 9436
rect 38192 9380 38240 9436
rect 38296 9380 38324 9436
rect 38004 7868 38324 9380
rect 38004 7812 38032 7868
rect 38088 7812 38136 7868
rect 38192 7812 38240 7868
rect 38296 7812 38324 7868
rect 38004 6300 38324 7812
rect 38004 6244 38032 6300
rect 38088 6244 38136 6300
rect 38192 6244 38240 6300
rect 38296 6244 38324 6300
rect 38004 4732 38324 6244
rect 38004 4676 38032 4732
rect 38088 4676 38136 4732
rect 38192 4676 38240 4732
rect 38296 4676 38324 4732
rect 19594 3076 19914 3892
rect 30492 3892 30548 3902
rect 30492 3556 30548 3836
rect 30492 3490 30548 3500
rect 38004 3164 38324 4676
rect 38004 3108 38032 3164
rect 38088 3108 38136 3164
rect 38192 3108 38240 3164
rect 38296 3108 38324 3164
rect 38004 3076 38324 3108
rect 56414 36876 56734 36908
rect 56414 36820 56442 36876
rect 56498 36820 56546 36876
rect 56602 36820 56650 36876
rect 56706 36820 56734 36876
rect 56414 35308 56734 36820
rect 56414 35252 56442 35308
rect 56498 35252 56546 35308
rect 56602 35252 56650 35308
rect 56706 35252 56734 35308
rect 56414 33740 56734 35252
rect 56414 33684 56442 33740
rect 56498 33684 56546 33740
rect 56602 33684 56650 33740
rect 56706 33684 56734 33740
rect 56414 32172 56734 33684
rect 56414 32116 56442 32172
rect 56498 32116 56546 32172
rect 56602 32116 56650 32172
rect 56706 32116 56734 32172
rect 56414 30604 56734 32116
rect 56414 30548 56442 30604
rect 56498 30548 56546 30604
rect 56602 30548 56650 30604
rect 56706 30548 56734 30604
rect 56414 29036 56734 30548
rect 56414 28980 56442 29036
rect 56498 28980 56546 29036
rect 56602 28980 56650 29036
rect 56706 28980 56734 29036
rect 56414 27468 56734 28980
rect 56414 27412 56442 27468
rect 56498 27412 56546 27468
rect 56602 27412 56650 27468
rect 56706 27412 56734 27468
rect 56414 25900 56734 27412
rect 56414 25844 56442 25900
rect 56498 25844 56546 25900
rect 56602 25844 56650 25900
rect 56706 25844 56734 25900
rect 56414 24332 56734 25844
rect 56414 24276 56442 24332
rect 56498 24276 56546 24332
rect 56602 24276 56650 24332
rect 56706 24276 56734 24332
rect 56414 22764 56734 24276
rect 56414 22708 56442 22764
rect 56498 22708 56546 22764
rect 56602 22708 56650 22764
rect 56706 22708 56734 22764
rect 56414 21196 56734 22708
rect 56414 21140 56442 21196
rect 56498 21140 56546 21196
rect 56602 21140 56650 21196
rect 56706 21140 56734 21196
rect 56414 19628 56734 21140
rect 56414 19572 56442 19628
rect 56498 19572 56546 19628
rect 56602 19572 56650 19628
rect 56706 19572 56734 19628
rect 56414 18060 56734 19572
rect 56414 18004 56442 18060
rect 56498 18004 56546 18060
rect 56602 18004 56650 18060
rect 56706 18004 56734 18060
rect 56414 16492 56734 18004
rect 56414 16436 56442 16492
rect 56498 16436 56546 16492
rect 56602 16436 56650 16492
rect 56706 16436 56734 16492
rect 56414 14924 56734 16436
rect 56414 14868 56442 14924
rect 56498 14868 56546 14924
rect 56602 14868 56650 14924
rect 56706 14868 56734 14924
rect 56414 13356 56734 14868
rect 56414 13300 56442 13356
rect 56498 13300 56546 13356
rect 56602 13300 56650 13356
rect 56706 13300 56734 13356
rect 56414 11788 56734 13300
rect 56414 11732 56442 11788
rect 56498 11732 56546 11788
rect 56602 11732 56650 11788
rect 56706 11732 56734 11788
rect 56414 10220 56734 11732
rect 56414 10164 56442 10220
rect 56498 10164 56546 10220
rect 56602 10164 56650 10220
rect 56706 10164 56734 10220
rect 56414 8652 56734 10164
rect 56414 8596 56442 8652
rect 56498 8596 56546 8652
rect 56602 8596 56650 8652
rect 56706 8596 56734 8652
rect 56414 7084 56734 8596
rect 56414 7028 56442 7084
rect 56498 7028 56546 7084
rect 56602 7028 56650 7084
rect 56706 7028 56734 7084
rect 56414 5516 56734 7028
rect 56414 5460 56442 5516
rect 56498 5460 56546 5516
rect 56602 5460 56650 5516
rect 56706 5460 56734 5516
rect 56414 3948 56734 5460
rect 56414 3892 56442 3948
rect 56498 3892 56546 3948
rect 56602 3892 56650 3948
rect 56706 3892 56734 3948
rect 56414 3076 56734 3892
rect 74824 36092 75144 36908
rect 74824 36036 74852 36092
rect 74908 36036 74956 36092
rect 75012 36036 75060 36092
rect 75116 36036 75144 36092
rect 74824 34524 75144 36036
rect 74824 34468 74852 34524
rect 74908 34468 74956 34524
rect 75012 34468 75060 34524
rect 75116 34468 75144 34524
rect 74824 32956 75144 34468
rect 74824 32900 74852 32956
rect 74908 32900 74956 32956
rect 75012 32900 75060 32956
rect 75116 32900 75144 32956
rect 74824 31388 75144 32900
rect 74824 31332 74852 31388
rect 74908 31332 74956 31388
rect 75012 31332 75060 31388
rect 75116 31332 75144 31388
rect 74824 29820 75144 31332
rect 74824 29764 74852 29820
rect 74908 29764 74956 29820
rect 75012 29764 75060 29820
rect 75116 29764 75144 29820
rect 74824 28252 75144 29764
rect 74824 28196 74852 28252
rect 74908 28196 74956 28252
rect 75012 28196 75060 28252
rect 75116 28196 75144 28252
rect 74824 26684 75144 28196
rect 74824 26628 74852 26684
rect 74908 26628 74956 26684
rect 75012 26628 75060 26684
rect 75116 26628 75144 26684
rect 74824 25116 75144 26628
rect 74824 25060 74852 25116
rect 74908 25060 74956 25116
rect 75012 25060 75060 25116
rect 75116 25060 75144 25116
rect 74824 23548 75144 25060
rect 74824 23492 74852 23548
rect 74908 23492 74956 23548
rect 75012 23492 75060 23548
rect 75116 23492 75144 23548
rect 74824 21980 75144 23492
rect 74824 21924 74852 21980
rect 74908 21924 74956 21980
rect 75012 21924 75060 21980
rect 75116 21924 75144 21980
rect 74824 20412 75144 21924
rect 74824 20356 74852 20412
rect 74908 20356 74956 20412
rect 75012 20356 75060 20412
rect 75116 20356 75144 20412
rect 74824 18844 75144 20356
rect 74824 18788 74852 18844
rect 74908 18788 74956 18844
rect 75012 18788 75060 18844
rect 75116 18788 75144 18844
rect 74824 17276 75144 18788
rect 74824 17220 74852 17276
rect 74908 17220 74956 17276
rect 75012 17220 75060 17276
rect 75116 17220 75144 17276
rect 74824 15708 75144 17220
rect 74824 15652 74852 15708
rect 74908 15652 74956 15708
rect 75012 15652 75060 15708
rect 75116 15652 75144 15708
rect 74824 14140 75144 15652
rect 74824 14084 74852 14140
rect 74908 14084 74956 14140
rect 75012 14084 75060 14140
rect 75116 14084 75144 14140
rect 74824 12572 75144 14084
rect 74824 12516 74852 12572
rect 74908 12516 74956 12572
rect 75012 12516 75060 12572
rect 75116 12516 75144 12572
rect 74824 11004 75144 12516
rect 74824 10948 74852 11004
rect 74908 10948 74956 11004
rect 75012 10948 75060 11004
rect 75116 10948 75144 11004
rect 74824 9436 75144 10948
rect 74824 9380 74852 9436
rect 74908 9380 74956 9436
rect 75012 9380 75060 9436
rect 75116 9380 75144 9436
rect 74824 7868 75144 9380
rect 74824 7812 74852 7868
rect 74908 7812 74956 7868
rect 75012 7812 75060 7868
rect 75116 7812 75144 7868
rect 74824 6300 75144 7812
rect 74824 6244 74852 6300
rect 74908 6244 74956 6300
rect 75012 6244 75060 6300
rect 75116 6244 75144 6300
rect 74824 4732 75144 6244
rect 93234 36876 93554 36908
rect 93234 36820 93262 36876
rect 93318 36820 93366 36876
rect 93422 36820 93470 36876
rect 93526 36820 93554 36876
rect 93234 35308 93554 36820
rect 93234 35252 93262 35308
rect 93318 35252 93366 35308
rect 93422 35252 93470 35308
rect 93526 35252 93554 35308
rect 93234 33740 93554 35252
rect 93234 33684 93262 33740
rect 93318 33684 93366 33740
rect 93422 33684 93470 33740
rect 93526 33684 93554 33740
rect 93234 32172 93554 33684
rect 93234 32116 93262 32172
rect 93318 32116 93366 32172
rect 93422 32116 93470 32172
rect 93526 32116 93554 32172
rect 93234 30604 93554 32116
rect 93234 30548 93262 30604
rect 93318 30548 93366 30604
rect 93422 30548 93470 30604
rect 93526 30548 93554 30604
rect 93234 29036 93554 30548
rect 93234 28980 93262 29036
rect 93318 28980 93366 29036
rect 93422 28980 93470 29036
rect 93526 28980 93554 29036
rect 93234 27468 93554 28980
rect 93234 27412 93262 27468
rect 93318 27412 93366 27468
rect 93422 27412 93470 27468
rect 93526 27412 93554 27468
rect 93234 25900 93554 27412
rect 93234 25844 93262 25900
rect 93318 25844 93366 25900
rect 93422 25844 93470 25900
rect 93526 25844 93554 25900
rect 93234 24332 93554 25844
rect 93234 24276 93262 24332
rect 93318 24276 93366 24332
rect 93422 24276 93470 24332
rect 93526 24276 93554 24332
rect 93234 22764 93554 24276
rect 93234 22708 93262 22764
rect 93318 22708 93366 22764
rect 93422 22708 93470 22764
rect 93526 22708 93554 22764
rect 93234 21196 93554 22708
rect 93234 21140 93262 21196
rect 93318 21140 93366 21196
rect 93422 21140 93470 21196
rect 93526 21140 93554 21196
rect 93234 19628 93554 21140
rect 93234 19572 93262 19628
rect 93318 19572 93366 19628
rect 93422 19572 93470 19628
rect 93526 19572 93554 19628
rect 93234 18060 93554 19572
rect 93234 18004 93262 18060
rect 93318 18004 93366 18060
rect 93422 18004 93470 18060
rect 93526 18004 93554 18060
rect 93234 16492 93554 18004
rect 93234 16436 93262 16492
rect 93318 16436 93366 16492
rect 93422 16436 93470 16492
rect 93526 16436 93554 16492
rect 93234 14924 93554 16436
rect 93234 14868 93262 14924
rect 93318 14868 93366 14924
rect 93422 14868 93470 14924
rect 93526 14868 93554 14924
rect 93234 13356 93554 14868
rect 93234 13300 93262 13356
rect 93318 13300 93366 13356
rect 93422 13300 93470 13356
rect 93526 13300 93554 13356
rect 93234 11788 93554 13300
rect 93234 11732 93262 11788
rect 93318 11732 93366 11788
rect 93422 11732 93470 11788
rect 93526 11732 93554 11788
rect 93234 10220 93554 11732
rect 93234 10164 93262 10220
rect 93318 10164 93366 10220
rect 93422 10164 93470 10220
rect 93526 10164 93554 10220
rect 93234 8652 93554 10164
rect 93234 8596 93262 8652
rect 93318 8596 93366 8652
rect 93422 8596 93470 8652
rect 93526 8596 93554 8652
rect 93234 7084 93554 8596
rect 93234 7028 93262 7084
rect 93318 7028 93366 7084
rect 93422 7028 93470 7084
rect 93526 7028 93554 7084
rect 88956 6020 89012 6030
rect 89012 5964 89460 6020
rect 88956 5954 89012 5964
rect 89404 5908 89460 5964
rect 89404 5842 89460 5852
rect 74824 4676 74852 4732
rect 74908 4676 74956 4732
rect 75012 4676 75060 4732
rect 75116 4676 75144 4732
rect 74824 3164 75144 4676
rect 74824 3108 74852 3164
rect 74908 3108 74956 3164
rect 75012 3108 75060 3164
rect 75116 3108 75144 3164
rect 74824 3076 75144 3108
rect 93234 5516 93554 7028
rect 93234 5460 93262 5516
rect 93318 5460 93366 5516
rect 93422 5460 93470 5516
rect 93526 5460 93554 5516
rect 93234 3948 93554 5460
rect 93234 3892 93262 3948
rect 93318 3892 93366 3948
rect 93422 3892 93470 3948
rect 93526 3892 93554 3948
rect 93234 3076 93554 3892
rect 111644 36092 111964 36908
rect 111644 36036 111672 36092
rect 111728 36036 111776 36092
rect 111832 36036 111880 36092
rect 111936 36036 111964 36092
rect 111644 34524 111964 36036
rect 111644 34468 111672 34524
rect 111728 34468 111776 34524
rect 111832 34468 111880 34524
rect 111936 34468 111964 34524
rect 111644 32956 111964 34468
rect 111644 32900 111672 32956
rect 111728 32900 111776 32956
rect 111832 32900 111880 32956
rect 111936 32900 111964 32956
rect 111644 31388 111964 32900
rect 111644 31332 111672 31388
rect 111728 31332 111776 31388
rect 111832 31332 111880 31388
rect 111936 31332 111964 31388
rect 111644 29820 111964 31332
rect 111644 29764 111672 29820
rect 111728 29764 111776 29820
rect 111832 29764 111880 29820
rect 111936 29764 111964 29820
rect 111644 28252 111964 29764
rect 111644 28196 111672 28252
rect 111728 28196 111776 28252
rect 111832 28196 111880 28252
rect 111936 28196 111964 28252
rect 111644 26684 111964 28196
rect 111644 26628 111672 26684
rect 111728 26628 111776 26684
rect 111832 26628 111880 26684
rect 111936 26628 111964 26684
rect 111644 25116 111964 26628
rect 111644 25060 111672 25116
rect 111728 25060 111776 25116
rect 111832 25060 111880 25116
rect 111936 25060 111964 25116
rect 111644 23548 111964 25060
rect 111644 23492 111672 23548
rect 111728 23492 111776 23548
rect 111832 23492 111880 23548
rect 111936 23492 111964 23548
rect 111644 21980 111964 23492
rect 111644 21924 111672 21980
rect 111728 21924 111776 21980
rect 111832 21924 111880 21980
rect 111936 21924 111964 21980
rect 111644 20412 111964 21924
rect 111644 20356 111672 20412
rect 111728 20356 111776 20412
rect 111832 20356 111880 20412
rect 111936 20356 111964 20412
rect 111644 18844 111964 20356
rect 111644 18788 111672 18844
rect 111728 18788 111776 18844
rect 111832 18788 111880 18844
rect 111936 18788 111964 18844
rect 111644 17276 111964 18788
rect 111644 17220 111672 17276
rect 111728 17220 111776 17276
rect 111832 17220 111880 17276
rect 111936 17220 111964 17276
rect 111644 15708 111964 17220
rect 111644 15652 111672 15708
rect 111728 15652 111776 15708
rect 111832 15652 111880 15708
rect 111936 15652 111964 15708
rect 111644 14140 111964 15652
rect 111644 14084 111672 14140
rect 111728 14084 111776 14140
rect 111832 14084 111880 14140
rect 111936 14084 111964 14140
rect 111644 12572 111964 14084
rect 111644 12516 111672 12572
rect 111728 12516 111776 12572
rect 111832 12516 111880 12572
rect 111936 12516 111964 12572
rect 111644 11004 111964 12516
rect 111644 10948 111672 11004
rect 111728 10948 111776 11004
rect 111832 10948 111880 11004
rect 111936 10948 111964 11004
rect 111644 9436 111964 10948
rect 111644 9380 111672 9436
rect 111728 9380 111776 9436
rect 111832 9380 111880 9436
rect 111936 9380 111964 9436
rect 111644 7868 111964 9380
rect 111644 7812 111672 7868
rect 111728 7812 111776 7868
rect 111832 7812 111880 7868
rect 111936 7812 111964 7868
rect 111644 6300 111964 7812
rect 111644 6244 111672 6300
rect 111728 6244 111776 6300
rect 111832 6244 111880 6300
rect 111936 6244 111964 6300
rect 111644 4732 111964 6244
rect 111644 4676 111672 4732
rect 111728 4676 111776 4732
rect 111832 4676 111880 4732
rect 111936 4676 111964 4732
rect 110908 3780 110964 3790
rect 111356 3780 111412 3790
rect 110964 3724 111356 3780
rect 110908 3714 110964 3724
rect 111356 3714 111412 3724
rect 111644 3164 111964 4676
rect 111644 3108 111672 3164
rect 111728 3108 111776 3164
rect 111832 3108 111880 3164
rect 111936 3108 111964 3164
rect 111644 3076 111964 3108
rect 130054 36876 130374 36908
rect 130054 36820 130082 36876
rect 130138 36820 130186 36876
rect 130242 36820 130290 36876
rect 130346 36820 130374 36876
rect 130054 35308 130374 36820
rect 130054 35252 130082 35308
rect 130138 35252 130186 35308
rect 130242 35252 130290 35308
rect 130346 35252 130374 35308
rect 130054 33740 130374 35252
rect 130054 33684 130082 33740
rect 130138 33684 130186 33740
rect 130242 33684 130290 33740
rect 130346 33684 130374 33740
rect 130054 32172 130374 33684
rect 130054 32116 130082 32172
rect 130138 32116 130186 32172
rect 130242 32116 130290 32172
rect 130346 32116 130374 32172
rect 130054 30604 130374 32116
rect 130054 30548 130082 30604
rect 130138 30548 130186 30604
rect 130242 30548 130290 30604
rect 130346 30548 130374 30604
rect 130054 29036 130374 30548
rect 130054 28980 130082 29036
rect 130138 28980 130186 29036
rect 130242 28980 130290 29036
rect 130346 28980 130374 29036
rect 130054 27468 130374 28980
rect 130054 27412 130082 27468
rect 130138 27412 130186 27468
rect 130242 27412 130290 27468
rect 130346 27412 130374 27468
rect 130054 25900 130374 27412
rect 130054 25844 130082 25900
rect 130138 25844 130186 25900
rect 130242 25844 130290 25900
rect 130346 25844 130374 25900
rect 130054 24332 130374 25844
rect 130054 24276 130082 24332
rect 130138 24276 130186 24332
rect 130242 24276 130290 24332
rect 130346 24276 130374 24332
rect 130054 22764 130374 24276
rect 130054 22708 130082 22764
rect 130138 22708 130186 22764
rect 130242 22708 130290 22764
rect 130346 22708 130374 22764
rect 130054 21196 130374 22708
rect 130054 21140 130082 21196
rect 130138 21140 130186 21196
rect 130242 21140 130290 21196
rect 130346 21140 130374 21196
rect 130054 19628 130374 21140
rect 130054 19572 130082 19628
rect 130138 19572 130186 19628
rect 130242 19572 130290 19628
rect 130346 19572 130374 19628
rect 130054 18060 130374 19572
rect 130054 18004 130082 18060
rect 130138 18004 130186 18060
rect 130242 18004 130290 18060
rect 130346 18004 130374 18060
rect 130054 16492 130374 18004
rect 130054 16436 130082 16492
rect 130138 16436 130186 16492
rect 130242 16436 130290 16492
rect 130346 16436 130374 16492
rect 130054 14924 130374 16436
rect 130054 14868 130082 14924
rect 130138 14868 130186 14924
rect 130242 14868 130290 14924
rect 130346 14868 130374 14924
rect 130054 13356 130374 14868
rect 130054 13300 130082 13356
rect 130138 13300 130186 13356
rect 130242 13300 130290 13356
rect 130346 13300 130374 13356
rect 130054 11788 130374 13300
rect 130054 11732 130082 11788
rect 130138 11732 130186 11788
rect 130242 11732 130290 11788
rect 130346 11732 130374 11788
rect 130054 10220 130374 11732
rect 130054 10164 130082 10220
rect 130138 10164 130186 10220
rect 130242 10164 130290 10220
rect 130346 10164 130374 10220
rect 130054 8652 130374 10164
rect 130054 8596 130082 8652
rect 130138 8596 130186 8652
rect 130242 8596 130290 8652
rect 130346 8596 130374 8652
rect 130054 7084 130374 8596
rect 130054 7028 130082 7084
rect 130138 7028 130186 7084
rect 130242 7028 130290 7084
rect 130346 7028 130374 7084
rect 130054 5516 130374 7028
rect 130054 5460 130082 5516
rect 130138 5460 130186 5516
rect 130242 5460 130290 5516
rect 130346 5460 130374 5516
rect 130054 3948 130374 5460
rect 130054 3892 130082 3948
rect 130138 3892 130186 3948
rect 130242 3892 130290 3948
rect 130346 3892 130374 3948
rect 148464 36092 148784 36908
rect 148464 36036 148492 36092
rect 148548 36036 148596 36092
rect 148652 36036 148700 36092
rect 148756 36036 148784 36092
rect 148464 34524 148784 36036
rect 148464 34468 148492 34524
rect 148548 34468 148596 34524
rect 148652 34468 148700 34524
rect 148756 34468 148784 34524
rect 148464 32956 148784 34468
rect 148464 32900 148492 32956
rect 148548 32900 148596 32956
rect 148652 32900 148700 32956
rect 148756 32900 148784 32956
rect 148464 31388 148784 32900
rect 148464 31332 148492 31388
rect 148548 31332 148596 31388
rect 148652 31332 148700 31388
rect 148756 31332 148784 31388
rect 148464 29820 148784 31332
rect 148464 29764 148492 29820
rect 148548 29764 148596 29820
rect 148652 29764 148700 29820
rect 148756 29764 148784 29820
rect 148464 28252 148784 29764
rect 148464 28196 148492 28252
rect 148548 28196 148596 28252
rect 148652 28196 148700 28252
rect 148756 28196 148784 28252
rect 148464 26684 148784 28196
rect 148464 26628 148492 26684
rect 148548 26628 148596 26684
rect 148652 26628 148700 26684
rect 148756 26628 148784 26684
rect 148464 25116 148784 26628
rect 148464 25060 148492 25116
rect 148548 25060 148596 25116
rect 148652 25060 148700 25116
rect 148756 25060 148784 25116
rect 148464 23548 148784 25060
rect 148464 23492 148492 23548
rect 148548 23492 148596 23548
rect 148652 23492 148700 23548
rect 148756 23492 148784 23548
rect 148464 21980 148784 23492
rect 148464 21924 148492 21980
rect 148548 21924 148596 21980
rect 148652 21924 148700 21980
rect 148756 21924 148784 21980
rect 148464 20412 148784 21924
rect 148464 20356 148492 20412
rect 148548 20356 148596 20412
rect 148652 20356 148700 20412
rect 148756 20356 148784 20412
rect 148464 18844 148784 20356
rect 148464 18788 148492 18844
rect 148548 18788 148596 18844
rect 148652 18788 148700 18844
rect 148756 18788 148784 18844
rect 148464 17276 148784 18788
rect 148464 17220 148492 17276
rect 148548 17220 148596 17276
rect 148652 17220 148700 17276
rect 148756 17220 148784 17276
rect 148464 15708 148784 17220
rect 148464 15652 148492 15708
rect 148548 15652 148596 15708
rect 148652 15652 148700 15708
rect 148756 15652 148784 15708
rect 148464 14140 148784 15652
rect 148464 14084 148492 14140
rect 148548 14084 148596 14140
rect 148652 14084 148700 14140
rect 148756 14084 148784 14140
rect 148464 12572 148784 14084
rect 148464 12516 148492 12572
rect 148548 12516 148596 12572
rect 148652 12516 148700 12572
rect 148756 12516 148784 12572
rect 148464 11004 148784 12516
rect 148464 10948 148492 11004
rect 148548 10948 148596 11004
rect 148652 10948 148700 11004
rect 148756 10948 148784 11004
rect 148464 9436 148784 10948
rect 148464 9380 148492 9436
rect 148548 9380 148596 9436
rect 148652 9380 148700 9436
rect 148756 9380 148784 9436
rect 148464 7868 148784 9380
rect 148464 7812 148492 7868
rect 148548 7812 148596 7868
rect 148652 7812 148700 7868
rect 148756 7812 148784 7868
rect 148464 6300 148784 7812
rect 148464 6244 148492 6300
rect 148548 6244 148596 6300
rect 148652 6244 148700 6300
rect 148756 6244 148784 6300
rect 148464 4732 148784 6244
rect 148464 4676 148492 4732
rect 148548 4676 148596 4732
rect 148652 4676 148700 4732
rect 148756 4676 148784 4732
rect 130054 3076 130374 3892
rect 130956 3892 131012 3902
rect 130956 3444 131012 3836
rect 130956 3378 131012 3388
rect 148464 3164 148784 4676
rect 148464 3108 148492 3164
rect 148548 3108 148596 3164
rect 148652 3108 148700 3164
rect 148756 3108 148784 3164
rect 148464 3076 148784 3108
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__042__I dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 131712 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__044__I0
timestamp 1669390400
transform -1 0 121520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__044__S
timestamp 1669390400
transform 1 0 123424 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__046__I0
timestamp 1669390400
transform 1 0 122080 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__046__S
timestamp 1669390400
transform -1 0 124432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__048__I0
timestamp 1669390400
transform 1 0 126784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__048__S
timestamp 1669390400
transform 1 0 126560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__050__I0
timestamp 1669390400
transform -1 0 126560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__050__S
timestamp 1669390400
transform -1 0 129360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__053__I0
timestamp 1669390400
transform -1 0 128352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__055__I0
timestamp 1669390400
transform -1 0 128912 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__057__I0
timestamp 1669390400
transform -1 0 130480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__059__I0
timestamp 1669390400
transform -1 0 132048 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__062__I0
timestamp 1669390400
transform -1 0 134064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__064__I0
timestamp 1669390400
transform -1 0 135968 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__066__I0
timestamp 1669390400
transform 1 0 139776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__068__I0
timestamp 1669390400
transform -1 0 141568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__I0
timestamp 1669390400
transform -1 0 140000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__071__S
timestamp 1669390400
transform 1 0 140336 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__073__I0
timestamp 1669390400
transform -1 0 137648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__073__S
timestamp 1669390400
transform 1 0 136976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__075__I0
timestamp 1669390400
transform 1 0 136192 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__075__S
timestamp 1669390400
transform -1 0 137872 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__I0
timestamp 1669390400
transform 1 0 106960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__I1
timestamp 1669390400
transform 1 0 105952 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__077__S
timestamp 1669390400
transform 1 0 107408 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__079__I
timestamp 1669390400
transform 1 0 129808 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__080__I
timestamp 1669390400
transform -1 0 103376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__I0
timestamp 1669390400
transform -1 0 94640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__081__S
timestamp 1669390400
transform 1 0 97104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__083__I0
timestamp 1669390400
transform 1 0 96432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__083__S
timestamp 1669390400
transform 1 0 99456 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__084__I
timestamp 1669390400
transform -1 0 100576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__I0
timestamp 1669390400
transform 1 0 96432 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__085__S
timestamp 1669390400
transform 1 0 99008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__087__I0
timestamp 1669390400
transform -1 0 98672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__087__S
timestamp 1669390400
transform 1 0 101024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__089__I
timestamp 1669390400
transform 1 0 109536 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__090__I0
timestamp 1669390400
transform -1 0 101584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__092__I0
timestamp 1669390400
transform 1 0 101920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__094__I0
timestamp 1669390400
transform -1 0 104496 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__096__I0
timestamp 1669390400
transform 1 0 107072 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__098__I
timestamp 1669390400
transform 1 0 111440 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__099__I0
timestamp 1669390400
transform -1 0 108864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__101__I0
timestamp 1669390400
transform 1 0 109088 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__102__I
timestamp 1669390400
transform 1 0 110656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__103__I0
timestamp 1669390400
transform 1 0 112224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__105__I0
timestamp 1669390400
transform -1 0 112784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__107__I
timestamp 1669390400
transform 1 0 120176 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__I0
timestamp 1669390400
transform -1 0 114800 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__110__I0
timestamp 1669390400
transform 1 0 115248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__I0
timestamp 1669390400
transform 1 0 115696 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__114__I0
timestamp 1669390400
transform -1 0 118048 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__116__I
timestamp 1669390400
transform -1 0 76608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__117__I
timestamp 1669390400
transform 1 0 78512 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__I
timestamp 1669390400
transform 1 0 80528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__I
timestamp 1669390400
transform 1 0 81424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__I
timestamp 1669390400
transform 1 0 83776 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__I
timestamp 1669390400
transform 1 0 86912 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__122__I
timestamp 1669390400
transform 1 0 86912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__I
timestamp 1669390400
transform 1 0 88144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__I
timestamp 1669390400
transform 1 0 89824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__125__I
timestamp 1669390400
transform 1 0 77616 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__126__I
timestamp 1669390400
transform 1 0 79408 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I
timestamp 1669390400
transform 1 0 82096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__I
timestamp 1669390400
transform -1 0 82880 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__I
timestamp 1669390400
transform -1 0 85456 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__130__I
timestamp 1669390400
transform 1 0 86016 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__131__I
timestamp 1669390400
transform 1 0 88368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__I
timestamp 1669390400
transform 1 0 90272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__133__I
timestamp 1669390400
transform 1 0 90720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__I
timestamp 1669390400
transform -1 0 72800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__I
timestamp 1669390400
transform 1 0 76160 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform 1 0 146832 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform -1 0 144368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform 1 0 146832 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1669390400
transform -1 0 147504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1669390400
transform 1 0 147280 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1669390400
transform -1 0 147056 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1669390400
transform -1 0 147056 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1669390400
transform 1 0 146832 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1669390400
transform -1 0 147056 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1669390400
transform 1 0 146832 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1669390400
transform 1 0 146832 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1669390400
transform -1 0 21840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1669390400
transform 1 0 40880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1669390400
transform 1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1669390400
transform -1 0 42000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1669390400
transform 1 0 45360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1669390400
transform -1 0 45584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1669390400
transform 1 0 48720 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1669390400
transform -1 0 48944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1669390400
transform 1 0 52640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1669390400
transform -1 0 52080 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1669390400
transform -1 0 53760 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1669390400
transform 1 0 25200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1669390400
transform 1 0 56896 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1669390400
transform -1 0 57344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1669390400
transform 1 0 60480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1669390400
transform -1 0 60480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1669390400
transform 1 0 64400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1669390400
transform -1 0 63840 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1669390400
transform -1 0 65520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1669390400
transform 1 0 68880 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1669390400
transform -1 0 69440 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1669390400
transform 1 0 71792 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1669390400
transform -1 0 25088 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1669390400
transform 1 0 72576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1669390400
transform 1 0 75712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1669390400
transform 1 0 29120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1669390400
transform 1 0 30240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1669390400
transform -1 0 30464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1669390400
transform 1 0 33040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1669390400
transform -1 0 33040 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1669390400
transform 1 0 36960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1669390400
transform -1 0 36960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1669390400
transform -1 0 92400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1669390400
transform 1 0 111776 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1669390400
transform 1 0 113456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1669390400
transform 1 0 113904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1669390400
transform -1 0 114912 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1669390400
transform -1 0 115472 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1669390400
transform 1 0 118496 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1669390400
transform 1 0 121520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1669390400
transform 1 0 121968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1669390400
transform -1 0 122752 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1669390400
transform -1 0 124320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1669390400
transform -1 0 94080 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1669390400
transform -1 0 126112 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1669390400
transform -1 0 127904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1669390400
transform 1 0 135296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1669390400
transform 1 0 134176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1669390400
transform 1 0 135744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1669390400
transform 1 0 136192 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1669390400
transform 1 0 136976 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1669390400
transform -1 0 139104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1669390400
transform 1 0 140896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1669390400
transform 1 0 141792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1669390400
transform -1 0 95312 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1669390400
transform 1 0 145040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1669390400
transform 1 0 146832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1669390400
transform 1 0 98000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1669390400
transform -1 0 99232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1669390400
transform -1 0 100800 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1669390400
transform -1 0 103152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1669390400
transform 1 0 106736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1669390400
transform 1 0 107856 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1669390400
transform 1 0 108192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output76_I
timestamp 1669390400
transform -1 0 8960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output77_I
timestamp 1669390400
transform -1 0 9856 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output78_I
timestamp 1669390400
transform -1 0 11424 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output79_I
timestamp 1669390400
transform 1 0 12992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output80_I
timestamp 1669390400
transform 1 0 15120 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output81_I
timestamp 1669390400
transform -1 0 17136 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output82_I
timestamp 1669390400
transform 1 0 18256 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output83_I
timestamp 1669390400
transform 1 0 20496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output84_I
timestamp 1669390400
transform -1 0 21504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output94_I
timestamp 1669390400
transform -1 0 6720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output96_I
timestamp 1669390400
transform 1 0 144368 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output97_I
timestamp 1669390400
transform 1 0 144368 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output98_I
timestamp 1669390400
transform -1 0 144368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output99_I
timestamp 1669390400
transform 1 0 144368 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output100_I
timestamp 1669390400
transform -1 0 144368 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output101_I
timestamp 1669390400
transform 1 0 144368 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output102_I
timestamp 1669390400
transform -1 0 144368 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output103_I
timestamp 1669390400
transform 1 0 144368 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output104_I
timestamp 1669390400
transform 1 0 144368 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output105_I
timestamp 1669390400
transform -1 0 144368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output106_I
timestamp 1669390400
transform 1 0 144368 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output107_I
timestamp 1669390400
transform -1 0 144368 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output108_I
timestamp 1669390400
transform -1 0 144368 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output109_I
timestamp 1669390400
transform 1 0 144368 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output110_I
timestamp 1669390400
transform -1 0 144368 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output111_I
timestamp 1669390400
transform 1 0 144368 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output112_I
timestamp 1669390400
transform 1 0 144368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output113_I
timestamp 1669390400
transform -1 0 144368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output114_I
timestamp 1669390400
transform 1 0 144368 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output115_I
timestamp 1669390400
transform -1 0 144368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output116_I
timestamp 1669390400
transform -1 0 143920 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output117_I
timestamp 1669390400
transform 1 0 147056 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output118_I
timestamp 1669390400
transform 1 0 144368 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output119_I
timestamp 1669390400
transform 1 0 142128 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output120_I
timestamp 1669390400
transform 1 0 146608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output121_I
timestamp 1669390400
transform 1 0 144368 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output122_I
timestamp 1669390400
transform -1 0 144368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output123_I
timestamp 1669390400
transform 1 0 144368 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output124_I
timestamp 1669390400
transform -1 0 144368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output125_I
timestamp 1669390400
transform 1 0 144368 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output126_I
timestamp 1669390400
transform -1 0 144368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output127_I
timestamp 1669390400
transform 1 0 144368 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1669390400
transform 1 0 5488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7168 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54
timestamp 1669390400
transform 1 0 7392 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_69
timestamp 1669390400
transform 1 0 9072 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72
timestamp 1669390400
transform 1 0 9408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88
timestamp 1669390400
transform 1 0 11200 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_107
timestamp 1669390400
transform 1 0 13328 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_123
timestamp 1669390400
transform 1 0 15120 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_157
timestamp 1669390400
transform 1 0 18928 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_159
timestamp 1669390400
transform 1 0 19152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_174
timestamp 1669390400
transform 1 0 20832 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1669390400
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_180 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 21504 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_188 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 22400 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_192
timestamp 1669390400
transform 1 0 22848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_215
timestamp 1669390400
transform 1 0 25424 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_223
timestamp 1669390400
transform 1 0 26320 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_227
timestamp 1669390400
transform 1 0 26768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_244
timestamp 1669390400
transform 1 0 28672 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_250
timestamp 1669390400
transform 1 0 29344 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_260
timestamp 1669390400
transform 1 0 30464 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_262
timestamp 1669390400
transform 1 0 30688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1669390400
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_285
timestamp 1669390400
transform 1 0 33264 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_293
timestamp 1669390400
transform 1 0 34160 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_297
timestamp 1669390400
transform 1 0 34608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1669390400
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_320
timestamp 1669390400
transform 1 0 37184 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_328
timestamp 1669390400
transform 1 0 38080 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_332
timestamp 1669390400
transform 1 0 38528 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1669390400
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_355
timestamp 1669390400
transform 1 0 41104 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_359
timestamp 1669390400
transform 1 0 41552 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_363
timestamp 1669390400
transform 1 0 42000 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_381
timestamp 1669390400
transform 1 0 44016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_391
timestamp 1669390400
transform 1 0 45136 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_395
timestamp 1669390400
transform 1 0 45584 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1669390400
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_422
timestamp 1669390400
transform 1 0 48608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_425
timestamp 1669390400
transform 1 0 48944 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_433
timestamp 1669390400
transform 1 0 49840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_437
timestamp 1669390400
transform 1 0 50288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_454
timestamp 1669390400
transform 1 0 52192 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_457
timestamp 1669390400
transform 1 0 52528 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_460
timestamp 1669390400
transform 1 0 52864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_464
timestamp 1669390400
transform 1 0 53312 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_468
timestamp 1669390400
transform 1 0 53760 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_486
timestamp 1669390400
transform 1 0 55776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_492
timestamp 1669390400
transform 1 0 56448 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_496
timestamp 1669390400
transform 1 0 56896 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_500
timestamp 1669390400
transform 1 0 57344 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_524
timestamp 1669390400
transform 1 0 60032 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_527
timestamp 1669390400
transform 1 0 60368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_530
timestamp 1669390400
transform 1 0 60704 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_538
timestamp 1669390400
transform 1 0 61600 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_542
timestamp 1669390400
transform 1 0 62048 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_559
timestamp 1669390400
transform 1 0 63952 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_562
timestamp 1669390400
transform 1 0 64288 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_565
timestamp 1669390400
transform 1 0 64624 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_569
timestamp 1669390400
transform 1 0 65072 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_573
timestamp 1669390400
transform 1 0 65520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_591
timestamp 1669390400
transform 1 0 67536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_597
timestamp 1669390400
transform 1 0 68208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_601
timestamp 1669390400
transform 1 0 68656 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_605
timestamp 1669390400
transform 1 0 69104 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_629
timestamp 1669390400
transform 1 0 71792 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_632
timestamp 1669390400
transform 1 0 72128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_638
timestamp 1669390400
transform 1 0 72800 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_646
timestamp 1669390400
transform 1 0 73696 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_664
timestamp 1669390400
transform 1 0 75712 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_667
timestamp 1669390400
transform 1 0 76048 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_682
timestamp 1669390400
transform 1 0 77728 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_698
timestamp 1669390400
transform 1 0 79520 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_702
timestamp 1669390400
transform 1 0 79968 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_717
timestamp 1669390400
transform 1 0 81648 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_733
timestamp 1669390400
transform 1 0 83440 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_737
timestamp 1669390400
transform 1 0 83888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_739
timestamp 1669390400
transform 1 0 84112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_754
timestamp 1669390400
transform 1 0 85792 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_762
timestamp 1669390400
transform 1 0 86688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_766
timestamp 1669390400
transform 1 0 87136 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_772
timestamp 1669390400
transform 1 0 87808 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_787
timestamp 1669390400
transform 1 0 89488 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_803
timestamp 1669390400
transform 1 0 91280 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_807
timestamp 1669390400
transform 1 0 91728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_813
timestamp 1669390400
transform 1 0 92400 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_831
timestamp 1669390400
transform 1 0 94416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_835
timestamp 1669390400
transform 1 0 94864 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_839
timestamp 1669390400
transform 1 0 95312 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_842
timestamp 1669390400
transform 1 0 95648 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_844
timestamp 1669390400
transform 1 0 95872 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_861
timestamp 1669390400
transform 1 0 97776 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_865
timestamp 1669390400
transform 1 0 98224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_869
timestamp 1669390400
transform 1 0 98672 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_871
timestamp 1669390400
transform 1 0 98896 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_874
timestamp 1669390400
transform 1 0 99232 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_877
timestamp 1669390400
transform 1 0 99568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_894
timestamp 1669390400
transform 1 0 101472 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_902
timestamp 1669390400
transform 1 0 102368 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_906
timestamp 1669390400
transform 1 0 102816 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_909
timestamp 1669390400
transform 1 0 103152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_912
timestamp 1669390400
transform 1 0 103488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_929
timestamp 1669390400
transform 1 0 105392 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_939
timestamp 1669390400
transform 1 0 106512 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_943
timestamp 1669390400
transform 1 0 106960 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_947
timestamp 1669390400
transform 1 0 107408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_964
timestamp 1669390400
transform 1 0 109312 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_968
timestamp 1669390400
transform 1 0 109760 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_978
timestamp 1669390400
transform 1 0 110880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_982
timestamp 1669390400
transform 1 0 111328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_999
timestamp 1669390400
transform 1 0 113232 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1003
timestamp 1669390400
transform 1 0 113680 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1007
timestamp 1669390400
transform 1 0 114128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1011
timestamp 1669390400
transform 1 0 114576 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1014
timestamp 1669390400
transform 1 0 114912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1017
timestamp 1669390400
transform 1 0 115248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1034
timestamp 1669390400
transform 1 0 117152 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1044
timestamp 1669390400
transform 1 0 118272 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1048
timestamp 1669390400
transform 1 0 118720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1052
timestamp 1669390400
transform 1 0 119168 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1054
timestamp 1669390400
transform 1 0 119392 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1071
timestamp 1669390400
transform 1 0 121296 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1075
timestamp 1669390400
transform 1 0 121744 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1079
timestamp 1669390400
transform 1 0 122192 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1081
timestamp 1669390400
transform 1 0 122416 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1084
timestamp 1669390400
transform 1 0 122752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1087
timestamp 1669390400
transform 1 0 123088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1104
timestamp 1669390400
transform 1 0 124992 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1114
timestamp 1669390400
transform 1 0 126112 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1118
timestamp 1669390400
transform 1 0 126560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1122
timestamp 1669390400
transform 1 0 127008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1139
timestamp 1669390400
transform 1 0 128912 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1143
timestamp 1669390400
transform 1 0 129360 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1145
timestamp 1669390400
transform 1 0 129584 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1154
timestamp 1669390400
transform 1 0 130592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1157
timestamp 1669390400
transform 1 0 130928 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1174
timestamp 1669390400
transform 1 0 132832 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1184
timestamp 1669390400
transform 1 0 133952 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1188
timestamp 1669390400
transform 1 0 134400 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1192
timestamp 1669390400
transform 1 0 134848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1209
timestamp 1669390400
transform 1 0 136752 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1213
timestamp 1669390400
transform 1 0 137200 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1217
timestamp 1669390400
transform 1 0 137648 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1224
timestamp 1669390400
transform 1 0 138432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1227
timestamp 1669390400
transform 1 0 138768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1244
timestamp 1669390400
transform 1 0 140672 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1248
timestamp 1669390400
transform 1 0 141120 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1252
timestamp 1669390400
transform 1 0 141568 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1256
timestamp 1669390400
transform 1 0 142016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1262
timestamp 1669390400
transform 1 0 142688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1264
timestamp 1669390400
transform 1 0 142912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1281
timestamp 1669390400
transform 1 0 144816 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1285
timestamp 1669390400
transform 1 0 145264 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1293
timestamp 1669390400
transform 1 0 146160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1297 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 146608 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_2
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_34
timestamp 1669390400
transform 1 0 5152 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_42
timestamp 1669390400
transform 1 0 6048 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_48
timestamp 1669390400
transform 1 0 6720 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_64
timestamp 1669390400
transform 1 0 8512 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_68
timestamp 1669390400
transform 1 0 8960 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_76
timestamp 1669390400
transform 1 0 9856 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_84
timestamp 1669390400
transform 1 0 10752 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_90
timestamp 1669390400
transform 1 0 11424 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_98
timestamp 1669390400
transform 1 0 12320 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_102
timestamp 1669390400
transform 1 0 12768 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_106
timestamp 1669390400
transform 1 0 13216 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_122
timestamp 1669390400
transform 1 0 15008 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_125
timestamp 1669390400
transform 1 0 15344 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_133
timestamp 1669390400
transform 1 0 16240 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_137
timestamp 1669390400
transform 1 0 16688 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1669390400
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_148
timestamp 1669390400
transform 1 0 17920 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_150
timestamp 1669390400
transform 1 0 18144 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_153
timestamp 1669390400
transform 1 0 18480 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_169
timestamp 1669390400
transform 1 0 20272 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_173
timestamp 1669390400
transform 1 0 20720 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_183
timestamp 1669390400
transform 1 0 21840 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_201
timestamp 1669390400
transform 1 0 23856 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_209
timestamp 1669390400
transform 1 0 24752 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1669390400
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_215
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_232
timestamp 1669390400
transform 1 0 27328 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_240
timestamp 1669390400
transform 1 0 28224 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_258
timestamp 1669390400
transform 1 0 30240 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_276
timestamp 1669390400
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_280
timestamp 1669390400
transform 1 0 32704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_306
timestamp 1669390400
transform 1 0 35616 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_314
timestamp 1669390400
transform 1 0 36512 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_318
timestamp 1669390400
transform 1 0 36960 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_336
timestamp 1669390400
transform 1 0 38976 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1669390400
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_374
timestamp 1669390400
transform 1 0 43232 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_376
timestamp 1669390400
transform 1 0 43456 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_393
timestamp 1669390400
transform 1 0 45360 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_411
timestamp 1669390400
transform 1 0 47376 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_419
timestamp 1669390400
transform 1 0 48272 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1669390400
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1669390400
transform 1 0 49280 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_445
timestamp 1669390400
transform 1 0 51184 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_449
timestamp 1669390400
transform 1 0 51632 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_453
timestamp 1669390400
transform 1 0 52080 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_471
timestamp 1669390400
transform 1 0 54096 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_479
timestamp 1669390400
transform 1 0 54992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_496
timestamp 1669390400
transform 1 0 56896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_499
timestamp 1669390400
transform 1 0 57232 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_516
timestamp 1669390400
transform 1 0 59136 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_524
timestamp 1669390400
transform 1 0 60032 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_528
timestamp 1669390400
transform 1 0 60480 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_546
timestamp 1669390400
transform 1 0 62496 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_562
timestamp 1669390400
transform 1 0 64288 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_566
timestamp 1669390400
transform 1 0 64736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_570
timestamp 1669390400
transform 1 0 65184 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_586
timestamp 1669390400
transform 1 0 66976 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_603
timestamp 1669390400
transform 1 0 68880 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_621
timestamp 1669390400
transform 1 0 70896 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_631
timestamp 1669390400
transform 1 0 72016 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_635
timestamp 1669390400
transform 1 0 72464 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_638
timestamp 1669390400
transform 1 0 72800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_641
timestamp 1669390400
transform 1 0 73136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_658
timestamp 1669390400
transform 1 0 75040 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_668
timestamp 1669390400
transform 1 0 76160 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_672
timestamp 1669390400
transform 1 0 76608 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_674
timestamp 1669390400
transform 1 0 76832 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_681
timestamp 1669390400
transform 1 0 77616 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_689
timestamp 1669390400
transform 1 0 78512 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_697
timestamp 1669390400
transform 1 0 79408 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_705
timestamp 1669390400
transform 1 0 80304 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_709
timestamp 1669390400
transform 1 0 80752 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_712
timestamp 1669390400
transform 1 0 81088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_719
timestamp 1669390400
transform 1 0 81872 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_723
timestamp 1669390400
transform 1 0 82320 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_739
timestamp 1669390400
transform 1 0 84112 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_747
timestamp 1669390400
transform 1 0 85008 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_751
timestamp 1669390400
transform 1 0 85456 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_769
timestamp 1669390400
transform 1 0 87472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_777
timestamp 1669390400
transform 1 0 88368 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_783
timestamp 1669390400
transform 1 0 89040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_790
timestamp 1669390400
transform 1 0 89824 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_798
timestamp 1669390400
transform 1 0 90720 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_814
timestamp 1669390400
transform 1 0 92512 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_822
timestamp 1669390400
transform 1 0 93408 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_828
timestamp 1669390400
transform 1 0 94080 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_846
timestamp 1669390400
transform 1 0 96096 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_848
timestamp 1669390400
transform 1 0 96320 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_851
timestamp 1669390400
transform 1 0 96656 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_854
timestamp 1669390400
transform 1 0 96992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_857
timestamp 1669390400
transform 1 0 97328 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_859
timestamp 1669390400
transform 1 0 97552 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_876
timestamp 1669390400
transform 1 0 99456 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_884
timestamp 1669390400
transform 1 0 100352 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_888
timestamp 1669390400
transform 1 0 100800 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_906
timestamp 1669390400
transform 1 0 102816 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_908
timestamp 1669390400
transform 1 0 103040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_911
timestamp 1669390400
transform 1 0 103376 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_921
timestamp 1669390400
transform 1 0 104496 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_925
timestamp 1669390400
transform 1 0 104944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_942
timestamp 1669390400
transform 1 0 106848 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_946
timestamp 1669390400
transform 1 0 107296 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_966
timestamp 1669390400
transform 1 0 109536 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_984
timestamp 1669390400
transform 1 0 111552 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_988
timestamp 1669390400
transform 1 0 112000 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_992
timestamp 1669390400
transform 1 0 112448 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_996
timestamp 1669390400
transform 1 0 112896 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1013
timestamp 1669390400
transform 1 0 114800 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1019
timestamp 1669390400
transform 1 0 115472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1023
timestamp 1669390400
transform 1 0 115920 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1041
timestamp 1669390400
transform 1 0 117936 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1059
timestamp 1669390400
transform 1 0 119952 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1063
timestamp 1669390400
transform 1 0 120400 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1067
timestamp 1669390400
transform 1 0 120848 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1069
timestamp 1669390400
transform 1 0 121072 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1086
timestamp 1669390400
transform 1 0 122976 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1092
timestamp 1669390400
transform 1 0 123648 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1098
timestamp 1669390400
transform 1 0 124320 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1116
timestamp 1669390400
transform 1 0 126336 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1133
timestamp 1669390400
transform 1 0 128240 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1135
timestamp 1669390400
transform 1 0 128464 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1138
timestamp 1669390400
transform 1 0 128800 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1155
timestamp 1669390400
transform 1 0 130704 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1159
timestamp 1669390400
transform 1 0 131152 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1176
timestamp 1669390400
transform 1 0 133056 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1194
timestamp 1669390400
transform 1 0 135072 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1198
timestamp 1669390400
transform 1 0 135520 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1202
timestamp 1669390400
transform 1 0 135968 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1206
timestamp 1669390400
transform 1 0 136416 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1209
timestamp 1669390400
transform 1 0 136752 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1226
timestamp 1669390400
transform 1 0 138656 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1230
timestamp 1669390400
transform 1 0 139104 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1234
timestamp 1669390400
transform 1 0 139552 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1251
timestamp 1669390400
transform 1 0 141456 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1269
timestamp 1669390400
transform 1 0 143472 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1277
timestamp 1669390400
transform 1 0 144368 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_1280
timestamp 1669390400
transform 1 0 144704 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_1297
timestamp 1669390400
transform 1 0 146608 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_1301
timestamp 1669390400
transform 1 0 147056 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_1309
timestamp 1669390400
transform 1 0 147952 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1669390400
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1669390400
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1669390400
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1669390400
transform 1 0 28560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_250
timestamp 1669390400
transform 1 0 29344 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_260
timestamp 1669390400
transform 1 0 30464 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_292
timestamp 1669390400
transform 1 0 34048 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_308
timestamp 1669390400
transform 1 0 35840 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_316
timestamp 1669390400
transform 1 0 36736 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_385
timestamp 1669390400
transform 1 0 44464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1669390400
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_395
timestamp 1669390400
transform 1 0 45584 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_459
timestamp 1669390400
transform 1 0 52752 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_463
timestamp 1669390400
transform 1 0 53200 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_495
timestamp 1669390400
transform 1 0 56784 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_498
timestamp 1669390400
transform 1 0 57120 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_530
timestamp 1669390400
transform 1 0 60704 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_534
timestamp 1669390400
transform 1 0 61152 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_550
timestamp 1669390400
transform 1 0 62944 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_554
timestamp 1669390400
transform 1 0 63392 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_558
timestamp 1669390400
transform 1 0 63840 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_576
timestamp 1669390400
transform 1 0 65856 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_592
timestamp 1669390400
transform 1 0 67648 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_600
timestamp 1669390400
transform 1 0 68544 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_602
timestamp 1669390400
transform 1 0 68768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_605
timestamp 1669390400
transform 1 0 69104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_608
timestamp 1669390400
transform 1 0 69440 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_640
timestamp 1669390400
transform 1 0 73024 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_656
timestamp 1669390400
transform 1 0 74816 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_666
timestamp 1669390400
transform 1 0 75936 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_670
timestamp 1669390400
transform 1 0 76384 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_676
timestamp 1669390400
transform 1 0 77056 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_680
timestamp 1669390400
transform 1 0 77504 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_683
timestamp 1669390400
transform 1 0 77840 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_687
timestamp 1669390400
transform 1 0 78288 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_691
timestamp 1669390400
transform 1 0 78736 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_695
timestamp 1669390400
transform 1 0 79184 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_699
timestamp 1669390400
transform 1 0 79632 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_713
timestamp 1669390400
transform 1 0 81200 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_717
timestamp 1669390400
transform 1 0 81648 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_719
timestamp 1669390400
transform 1 0 81872 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_726
timestamp 1669390400
transform 1 0 82656 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_734
timestamp 1669390400
transform 1 0 83552 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_738
timestamp 1669390400
transform 1 0 84000 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_742
timestamp 1669390400
transform 1 0 84448 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_744
timestamp 1669390400
transform 1 0 84672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_747
timestamp 1669390400
transform 1 0 85008 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_749
timestamp 1669390400
transform 1 0 85232 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_756
timestamp 1669390400
transform 1 0 86016 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_764
timestamp 1669390400
transform 1 0 86912 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_766
timestamp 1669390400
transform 1 0 87136 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_773
timestamp 1669390400
transform 1 0 87920 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_777
timestamp 1669390400
transform 1 0 88368 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_781
timestamp 1669390400
transform 1 0 88816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_788
timestamp 1669390400
transform 1 0 89600 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_792
timestamp 1669390400
transform 1 0 90048 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_796
timestamp 1669390400
transform 1 0 90496 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_800
timestamp 1669390400
transform 1 0 90944 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_818
timestamp 1669390400
transform 1 0 92960 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_826
timestamp 1669390400
transform 1 0 93856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_830
timestamp 1669390400
transform 1 0 94304 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_833
timestamp 1669390400
transform 1 0 94640 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_850
timestamp 1669390400
transform 1 0 96544 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_867
timestamp 1669390400
transform 1 0 98448 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_884
timestamp 1669390400
transform 1 0 100352 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_886
timestamp 1669390400
transform 1 0 100576 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_889
timestamp 1669390400
transform 1 0 100912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_892
timestamp 1669390400
transform 1 0 101248 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_894
timestamp 1669390400
transform 1 0 101472 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_910
timestamp 1669390400
transform 1 0 103264 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_927
timestamp 1669390400
transform 1 0 105168 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_944
timestamp 1669390400
transform 1 0 107072 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_952
timestamp 1669390400
transform 1 0 107968 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_956
timestamp 1669390400
transform 1 0 108416 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_960
timestamp 1669390400
transform 1 0 108864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_976
timestamp 1669390400
transform 1 0 110656 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_993
timestamp 1669390400
transform 1 0 112560 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1010
timestamp 1669390400
transform 1 0 114464 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1012
timestamp 1669390400
transform 1 0 114688 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1028
timestamp 1669390400
transform 1 0 116480 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1031
timestamp 1669390400
transform 1 0 116816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1047
timestamp 1669390400
transform 1 0 118608 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1055
timestamp 1669390400
transform 1 0 119504 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1063
timestamp 1669390400
transform 1 0 120400 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1073
timestamp 1669390400
transform 1 0 121520 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1090
timestamp 1669390400
transform 1 0 123424 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1098
timestamp 1669390400
transform 1 0 124320 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1102
timestamp 1669390400
transform 1 0 124768 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1118
timestamp 1669390400
transform 1 0 126560 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1122
timestamp 1669390400
transform 1 0 127008 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1132
timestamp 1669390400
transform 1 0 128128 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1149
timestamp 1669390400
transform 1 0 130032 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1151
timestamp 1669390400
transform 1 0 130256 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1167
timestamp 1669390400
transform 1 0 132048 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1173
timestamp 1669390400
transform 1 0 132720 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1182
timestamp 1669390400
transform 1 0 133728 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1184
timestamp 1669390400
transform 1 0 133952 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1200
timestamp 1669390400
transform 1 0 135744 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1217
timestamp 1669390400
transform 1 0 137648 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1234
timestamp 1669390400
transform 1 0 139552 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_1238
timestamp 1669390400
transform 1 0 140000 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1244
timestamp 1669390400
transform 1 0 140672 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1260
timestamp 1669390400
transform 1 0 142464 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_1262
timestamp 1669390400
transform 1 0 142688 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1279
timestamp 1669390400
transform 1 0 144592 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1297
timestamp 1669390400
transform 1 0 146608 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_1301
timestamp 1669390400
transform 1 0 147056 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_1305
timestamp 1669390400
transform 1 0 147504 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1669390400
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1669390400
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1669390400
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1669390400
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1669390400
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1669390400
transform 1 0 40544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1669390400
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_421
timestamp 1669390400
transform 1 0 48496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1669390400
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_428
timestamp 1669390400
transform 1 0 49280 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_492
timestamp 1669390400
transform 1 0 56448 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_496
timestamp 1669390400
transform 1 0 56896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_499
timestamp 1669390400
transform 1 0 57232 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_563
timestamp 1669390400
transform 1 0 64400 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_567
timestamp 1669390400
transform 1 0 64848 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_570
timestamp 1669390400
transform 1 0 65184 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_634
timestamp 1669390400
transform 1 0 72352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_638
timestamp 1669390400
transform 1 0 72800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_641
timestamp 1669390400
transform 1 0 73136 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_657
timestamp 1669390400
transform 1 0 74928 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_661
timestamp 1669390400
transform 1 0 75376 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_663
timestamp 1669390400
transform 1 0 75600 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_666
timestamp 1669390400
transform 1 0 75936 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_698
timestamp 1669390400
transform 1 0 79520 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_706
timestamp 1669390400
transform 1 0 80416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_712
timestamp 1669390400
transform 1 0 81088 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_720
timestamp 1669390400
transform 1 0 81984 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_724
timestamp 1669390400
transform 1 0 82432 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_728
timestamp 1669390400
transform 1 0 82880 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_744
timestamp 1669390400
transform 1 0 84672 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_752
timestamp 1669390400
transform 1 0 85568 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_758
timestamp 1669390400
transform 1 0 86240 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_762
timestamp 1669390400
transform 1 0 86688 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_766
timestamp 1669390400
transform 1 0 87136 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_774
timestamp 1669390400
transform 1 0 88032 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_776
timestamp 1669390400
transform 1 0 88256 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_779
timestamp 1669390400
transform 1 0 88592 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_783
timestamp 1669390400
transform 1 0 89040 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_847
timestamp 1669390400
transform 1 0 96208 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_851
timestamp 1669390400
transform 1 0 96656 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_854
timestamp 1669390400
transform 1 0 96992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_870
timestamp 1669390400
transform 1 0 98784 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_874
timestamp 1669390400
transform 1 0 99232 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_878
timestamp 1669390400
transform 1 0 99680 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_886
timestamp 1669390400
transform 1 0 100576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_890
timestamp 1669390400
transform 1 0 101024 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_892
timestamp 1669390400
transform 1 0 101248 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_895
timestamp 1669390400
transform 1 0 101584 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_897
timestamp 1669390400
transform 1 0 101808 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_900
timestamp 1669390400
transform 1 0 102144 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_917
timestamp 1669390400
transform 1 0 104048 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_921
timestamp 1669390400
transform 1 0 104496 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_925
timestamp 1669390400
transform 1 0 104944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_941
timestamp 1669390400
transform 1 0 106736 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_945
timestamp 1669390400
transform 1 0 107184 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_949
timestamp 1669390400
transform 1 0 107632 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_953
timestamp 1669390400
transform 1 0 108080 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_957
timestamp 1669390400
transform 1 0 108528 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_960
timestamp 1669390400
transform 1 0 108864 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_964
timestamp 1669390400
transform 1 0 109312 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_981
timestamp 1669390400
transform 1 0 111216 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_983
timestamp 1669390400
transform 1 0 111440 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_990
timestamp 1669390400
transform 1 0 112224 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_996
timestamp 1669390400
transform 1 0 112896 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1003
timestamp 1669390400
transform 1 0 113680 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1013
timestamp 1669390400
transform 1 0 114800 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1019
timestamp 1669390400
transform 1 0 115472 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1036
timestamp 1669390400
transform 1 0 117376 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1038
timestamp 1669390400
transform 1 0 117600 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1054
timestamp 1669390400
transform 1 0 119392 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1062
timestamp 1669390400
transform 1 0 120288 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1064
timestamp 1669390400
transform 1 0 120512 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1067
timestamp 1669390400
transform 1 0 120848 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1075
timestamp 1669390400
transform 1 0 121744 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1077
timestamp 1669390400
transform 1 0 121968 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1080
timestamp 1669390400
transform 1 0 122304 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1097
timestamp 1669390400
transform 1 0 124208 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1105
timestamp 1669390400
transform 1 0 125104 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1115
timestamp 1669390400
transform 1 0 126224 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1117
timestamp 1669390400
transform 1 0 126448 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1120
timestamp 1669390400
transform 1 0 126784 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1130
timestamp 1669390400
transform 1 0 127904 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1134
timestamp 1669390400
transform 1 0 128352 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1138
timestamp 1669390400
transform 1 0 128800 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1140
timestamp 1669390400
transform 1 0 129024 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1156
timestamp 1669390400
transform 1 0 130816 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1175
timestamp 1669390400
transform 1 0 132944 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1185
timestamp 1669390400
transform 1 0 134064 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_1193
timestamp 1669390400
transform 1 0 134960 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1197
timestamp 1669390400
transform 1 0 135408 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1199
timestamp 1669390400
transform 1 0 135632 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1202
timestamp 1669390400
transform 1 0 135968 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1206
timestamp 1669390400
transform 1 0 136416 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1209
timestamp 1669390400
transform 1 0 136752 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1216
timestamp 1669390400
transform 1 0 137536 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1218
timestamp 1669390400
transform 1 0 137760 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1234
timestamp 1669390400
transform 1 0 139552 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1251
timestamp 1669390400
transform 1 0 141456 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1259
timestamp 1669390400
transform 1 0 142352 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1277
timestamp 1669390400
transform 1 0 144368 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_1280
timestamp 1669390400
transform 1 0 144704 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1297
timestamp 1669390400
transform 1 0 146608 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_1301
timestamp 1669390400
transform 1 0 147056 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_1305
timestamp 1669390400
transform 1 0 147504 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1669390400
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1669390400
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1669390400
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1669390400
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1669390400
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1669390400
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1669390400
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1669390400
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_456
timestamp 1669390400
transform 1 0 52416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_460
timestamp 1669390400
transform 1 0 52864 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_463
timestamp 1669390400
transform 1 0 53200 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_527
timestamp 1669390400
transform 1 0 60368 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_531
timestamp 1669390400
transform 1 0 60816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_534
timestamp 1669390400
transform 1 0 61152 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_598
timestamp 1669390400
transform 1 0 68320 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_602
timestamp 1669390400
transform 1 0 68768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_605
timestamp 1669390400
transform 1 0 69104 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_669
timestamp 1669390400
transform 1 0 76272 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_673
timestamp 1669390400
transform 1 0 76720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_676
timestamp 1669390400
transform 1 0 77056 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_740
timestamp 1669390400
transform 1 0 84224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_744
timestamp 1669390400
transform 1 0 84672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_747
timestamp 1669390400
transform 1 0 85008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_811
timestamp 1669390400
transform 1 0 92176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_815
timestamp 1669390400
transform 1 0 92624 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_818
timestamp 1669390400
transform 1 0 92960 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_882
timestamp 1669390400
transform 1 0 100128 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_886
timestamp 1669390400
transform 1 0 100576 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_889
timestamp 1669390400
transform 1 0 100912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_896
timestamp 1669390400
transform 1 0 101696 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_904
timestamp 1669390400
transform 1 0 102592 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_908
timestamp 1669390400
transform 1 0 103040 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_915
timestamp 1669390400
transform 1 0 103824 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_923
timestamp 1669390400
transform 1 0 104720 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_925
timestamp 1669390400
transform 1 0 104944 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_932
timestamp 1669390400
transform 1 0 105728 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_936
timestamp 1669390400
transform 1 0 106176 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_952
timestamp 1669390400
transform 1 0 107968 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_956
timestamp 1669390400
transform 1 0 108416 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_960
timestamp 1669390400
transform 1 0 108864 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_968
timestamp 1669390400
transform 1 0 109760 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_972
timestamp 1669390400
transform 1 0 110208 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_981
timestamp 1669390400
transform 1 0 111216 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_985
timestamp 1669390400
transform 1 0 111664 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_995
timestamp 1669390400
transform 1 0 112784 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1027
timestamp 1669390400
transform 1 0 116368 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1031
timestamp 1669390400
transform 1 0 116816 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1038
timestamp 1669390400
transform 1 0 117600 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_1042
timestamp 1669390400
transform 1 0 118048 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_1074
timestamp 1669390400
transform 1 0 121632 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1090
timestamp 1669390400
transform 1 0 123424 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1094
timestamp 1669390400
transform 1 0 123872 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1096
timestamp 1669390400
transform 1 0 124096 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1099
timestamp 1669390400
transform 1 0 124432 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_1102
timestamp 1669390400
transform 1 0 124768 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1134
timestamp 1669390400
transform 1 0 128352 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1136
timestamp 1669390400
transform 1 0 128576 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1139
timestamp 1669390400
transform 1 0 128912 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1147
timestamp 1669390400
transform 1 0 129808 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1155
timestamp 1669390400
transform 1 0 130704 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1163
timestamp 1669390400
transform 1 0 131600 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1167
timestamp 1669390400
transform 1 0 132048 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1173
timestamp 1669390400
transform 1 0 132720 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1180
timestamp 1669390400
transform 1 0 133504 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1182
timestamp 1669390400
transform 1 0 133728 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_1185
timestamp 1669390400
transform 1 0 134064 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1201
timestamp 1669390400
transform 1 0 135856 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1209
timestamp 1669390400
transform 1 0 136752 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1213
timestamp 1669390400
transform 1 0 137200 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1217
timestamp 1669390400
transform 1 0 137648 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1234
timestamp 1669390400
transform 1 0 139552 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1238
timestamp 1669390400
transform 1 0 140000 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_1244
timestamp 1669390400
transform 1 0 140672 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1251
timestamp 1669390400
transform 1 0 141456 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1259
timestamp 1669390400
transform 1 0 142352 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1279
timestamp 1669390400
transform 1 0 144592 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_1297
timestamp 1669390400
transform 1 0 146608 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_4_1301
timestamp 1669390400
transform 1 0 147056 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_1309
timestamp 1669390400
transform 1 0 147952 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_66
timestamp 1669390400
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1669390400
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1669390400
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1669390400
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1669390400
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1669390400
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1669390400
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1669390400
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_421
timestamp 1669390400
transform 1 0 48496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1669390400
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_428
timestamp 1669390400
transform 1 0 49280 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_492
timestamp 1669390400
transform 1 0 56448 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1669390400
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_499
timestamp 1669390400
transform 1 0 57232 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_563
timestamp 1669390400
transform 1 0 64400 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_567
timestamp 1669390400
transform 1 0 64848 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_570
timestamp 1669390400
transform 1 0 65184 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_634
timestamp 1669390400
transform 1 0 72352 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_638
timestamp 1669390400
transform 1 0 72800 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_641
timestamp 1669390400
transform 1 0 73136 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_705
timestamp 1669390400
transform 1 0 80304 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_709
timestamp 1669390400
transform 1 0 80752 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_712
timestamp 1669390400
transform 1 0 81088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_776
timestamp 1669390400
transform 1 0 88256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_780
timestamp 1669390400
transform 1 0 88704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_783
timestamp 1669390400
transform 1 0 89040 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_847
timestamp 1669390400
transform 1 0 96208 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_851
timestamp 1669390400
transform 1 0 96656 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_854
timestamp 1669390400
transform 1 0 96992 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_918
timestamp 1669390400
transform 1 0 104160 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_922
timestamp 1669390400
transform 1 0 104608 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_925
timestamp 1669390400
transform 1 0 104944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_932
timestamp 1669390400
transform 1 0 105728 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_964
timestamp 1669390400
transform 1 0 109312 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_980
timestamp 1669390400
transform 1 0 111104 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_988
timestamp 1669390400
transform 1 0 112000 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_992
timestamp 1669390400
transform 1 0 112448 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_996
timestamp 1669390400
transform 1 0 112896 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1060
timestamp 1669390400
transform 1 0 120064 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1064
timestamp 1669390400
transform 1 0 120512 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_1067
timestamp 1669390400
transform 1 0 120848 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1131
timestamp 1669390400
transform 1 0 128016 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1135
timestamp 1669390400
transform 1 0 128464 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1138
timestamp 1669390400
transform 1 0 128800 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1146
timestamp 1669390400
transform 1 0 129696 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1149
timestamp 1669390400
transform 1 0 130032 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1153
timestamp 1669390400
transform 1 0 130480 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1155
timestamp 1669390400
transform 1 0 130704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1162
timestamp 1669390400
transform 1 0 131488 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_1166
timestamp 1669390400
transform 1 0 131936 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1198
timestamp 1669390400
transform 1 0 135520 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1206
timestamp 1669390400
transform 1 0 136416 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1209
timestamp 1669390400
transform 1 0 136752 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1219
timestamp 1669390400
transform 1 0 137872 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1223
timestamp 1669390400
transform 1 0 138320 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1231
timestamp 1669390400
transform 1 0 139216 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1239
timestamp 1669390400
transform 1 0 140112 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_1243
timestamp 1669390400
transform 1 0 140560 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1277
timestamp 1669390400
transform 1 0 144368 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_1280
timestamp 1669390400
transform 1 0 144704 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_1297
timestamp 1669390400
transform 1 0 146608 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_1301
timestamp 1669390400
transform 1 0 147056 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_1309
timestamp 1669390400
transform 1 0 147952 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1669390400
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1669390400
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1669390400
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1669390400
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1669390400
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1669390400
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1669390400
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_456
timestamp 1669390400
transform 1 0 52416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_460
timestamp 1669390400
transform 1 0 52864 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_463
timestamp 1669390400
transform 1 0 53200 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_527
timestamp 1669390400
transform 1 0 60368 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_531
timestamp 1669390400
transform 1 0 60816 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_534
timestamp 1669390400
transform 1 0 61152 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_598
timestamp 1669390400
transform 1 0 68320 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_602
timestamp 1669390400
transform 1 0 68768 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_605
timestamp 1669390400
transform 1 0 69104 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_669
timestamp 1669390400
transform 1 0 76272 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_673
timestamp 1669390400
transform 1 0 76720 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_676
timestamp 1669390400
transform 1 0 77056 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_740
timestamp 1669390400
transform 1 0 84224 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_744
timestamp 1669390400
transform 1 0 84672 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_747
timestamp 1669390400
transform 1 0 85008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_811
timestamp 1669390400
transform 1 0 92176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_815
timestamp 1669390400
transform 1 0 92624 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_818
timestamp 1669390400
transform 1 0 92960 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_882
timestamp 1669390400
transform 1 0 100128 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_886
timestamp 1669390400
transform 1 0 100576 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_889
timestamp 1669390400
transform 1 0 100912 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_953
timestamp 1669390400
transform 1 0 108080 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_957
timestamp 1669390400
transform 1 0 108528 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_960
timestamp 1669390400
transform 1 0 108864 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1024
timestamp 1669390400
transform 1 0 116032 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1028
timestamp 1669390400
transform 1 0 116480 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1031
timestamp 1669390400
transform 1 0 116816 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1095
timestamp 1669390400
transform 1 0 123984 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1099
timestamp 1669390400
transform 1 0 124432 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1102
timestamp 1669390400
transform 1 0 124768 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1166
timestamp 1669390400
transform 1 0 131936 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1170
timestamp 1669390400
transform 1 0 132384 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_1173
timestamp 1669390400
transform 1 0 132720 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1237
timestamp 1669390400
transform 1 0 139888 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1241
timestamp 1669390400
transform 1 0 140336 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_1244
timestamp 1669390400
transform 1 0 140672 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1276
timestamp 1669390400
transform 1 0 144256 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_1280
timestamp 1669390400
transform 1 0 144704 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_1297
timestamp 1669390400
transform 1 0 146608 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_1301
timestamp 1669390400
transform 1 0 147056 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_1309
timestamp 1669390400
transform 1 0 147952 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_66
timestamp 1669390400
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1669390400
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1669390400
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1669390400
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1669390400
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1669390400
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1669390400
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_421
timestamp 1669390400
transform 1 0 48496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_425
timestamp 1669390400
transform 1 0 48944 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_428
timestamp 1669390400
transform 1 0 49280 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_492
timestamp 1669390400
transform 1 0 56448 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1669390400
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_499
timestamp 1669390400
transform 1 0 57232 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_563
timestamp 1669390400
transform 1 0 64400 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_567
timestamp 1669390400
transform 1 0 64848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_570
timestamp 1669390400
transform 1 0 65184 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_634
timestamp 1669390400
transform 1 0 72352 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_638
timestamp 1669390400
transform 1 0 72800 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_641
timestamp 1669390400
transform 1 0 73136 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_705
timestamp 1669390400
transform 1 0 80304 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_709
timestamp 1669390400
transform 1 0 80752 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_712
timestamp 1669390400
transform 1 0 81088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_776
timestamp 1669390400
transform 1 0 88256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_780
timestamp 1669390400
transform 1 0 88704 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_783
timestamp 1669390400
transform 1 0 89040 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_847
timestamp 1669390400
transform 1 0 96208 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_851
timestamp 1669390400
transform 1 0 96656 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_854
timestamp 1669390400
transform 1 0 96992 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_918
timestamp 1669390400
transform 1 0 104160 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_922
timestamp 1669390400
transform 1 0 104608 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_925
timestamp 1669390400
transform 1 0 104944 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_989
timestamp 1669390400
transform 1 0 112112 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_993
timestamp 1669390400
transform 1 0 112560 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_996
timestamp 1669390400
transform 1 0 112896 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1060
timestamp 1669390400
transform 1 0 120064 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1064
timestamp 1669390400
transform 1 0 120512 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1067
timestamp 1669390400
transform 1 0 120848 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1131
timestamp 1669390400
transform 1 0 128016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1135
timestamp 1669390400
transform 1 0 128464 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1138
timestamp 1669390400
transform 1 0 128800 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1202
timestamp 1669390400
transform 1 0 135968 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1206
timestamp 1669390400
transform 1 0 136416 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_1209
timestamp 1669390400
transform 1 0 136752 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1273
timestamp 1669390400
transform 1 0 143920 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1277
timestamp 1669390400
transform 1 0 144368 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_1280
timestamp 1669390400
transform 1 0 144704 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_1297
timestamp 1669390400
transform 1 0 146608 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_1301
timestamp 1669390400
transform 1 0 147056 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_1309
timestamp 1669390400
transform 1 0 147952 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_101
timestamp 1669390400
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1669390400
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1669390400
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1669390400
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1669390400
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1669390400
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1669390400
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1669390400
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_456
timestamp 1669390400
transform 1 0 52416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1669390400
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_463
timestamp 1669390400
transform 1 0 53200 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_527
timestamp 1669390400
transform 1 0 60368 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_531
timestamp 1669390400
transform 1 0 60816 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_534
timestamp 1669390400
transform 1 0 61152 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_598
timestamp 1669390400
transform 1 0 68320 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_602
timestamp 1669390400
transform 1 0 68768 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_605
timestamp 1669390400
transform 1 0 69104 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_669
timestamp 1669390400
transform 1 0 76272 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_673
timestamp 1669390400
transform 1 0 76720 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_676
timestamp 1669390400
transform 1 0 77056 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_740
timestamp 1669390400
transform 1 0 84224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_744
timestamp 1669390400
transform 1 0 84672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_747
timestamp 1669390400
transform 1 0 85008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_811
timestamp 1669390400
transform 1 0 92176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_815
timestamp 1669390400
transform 1 0 92624 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_818
timestamp 1669390400
transform 1 0 92960 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_882
timestamp 1669390400
transform 1 0 100128 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_886
timestamp 1669390400
transform 1 0 100576 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_889
timestamp 1669390400
transform 1 0 100912 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_953
timestamp 1669390400
transform 1 0 108080 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_957
timestamp 1669390400
transform 1 0 108528 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_960
timestamp 1669390400
transform 1 0 108864 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1024
timestamp 1669390400
transform 1 0 116032 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1028
timestamp 1669390400
transform 1 0 116480 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1031
timestamp 1669390400
transform 1 0 116816 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1095
timestamp 1669390400
transform 1 0 123984 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1099
timestamp 1669390400
transform 1 0 124432 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1102
timestamp 1669390400
transform 1 0 124768 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1166
timestamp 1669390400
transform 1 0 131936 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1170
timestamp 1669390400
transform 1 0 132384 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_1173
timestamp 1669390400
transform 1 0 132720 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1237
timestamp 1669390400
transform 1 0 139888 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1241
timestamp 1669390400
transform 1 0 140336 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_1244
timestamp 1669390400
transform 1 0 140672 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1276
timestamp 1669390400
transform 1 0 144256 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_1280
timestamp 1669390400
transform 1 0 144704 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_1297
timestamp 1669390400
transform 1 0 146608 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_1301
timestamp 1669390400
transform 1 0 147056 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_1309
timestamp 1669390400
transform 1 0 147952 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_66
timestamp 1669390400
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1669390400
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1669390400
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1669390400
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1669390400
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1669390400
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1669390400
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_421
timestamp 1669390400
transform 1 0 48496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_425
timestamp 1669390400
transform 1 0 48944 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_428
timestamp 1669390400
transform 1 0 49280 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_492
timestamp 1669390400
transform 1 0 56448 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1669390400
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_499
timestamp 1669390400
transform 1 0 57232 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_563
timestamp 1669390400
transform 1 0 64400 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_567
timestamp 1669390400
transform 1 0 64848 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_570
timestamp 1669390400
transform 1 0 65184 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_634
timestamp 1669390400
transform 1 0 72352 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_638
timestamp 1669390400
transform 1 0 72800 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_641
timestamp 1669390400
transform 1 0 73136 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_705
timestamp 1669390400
transform 1 0 80304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_709
timestamp 1669390400
transform 1 0 80752 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_712
timestamp 1669390400
transform 1 0 81088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_776
timestamp 1669390400
transform 1 0 88256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_780
timestamp 1669390400
transform 1 0 88704 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_783
timestamp 1669390400
transform 1 0 89040 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_847
timestamp 1669390400
transform 1 0 96208 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_851
timestamp 1669390400
transform 1 0 96656 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_854
timestamp 1669390400
transform 1 0 96992 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_918
timestamp 1669390400
transform 1 0 104160 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_922
timestamp 1669390400
transform 1 0 104608 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_925
timestamp 1669390400
transform 1 0 104944 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_989
timestamp 1669390400
transform 1 0 112112 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_993
timestamp 1669390400
transform 1 0 112560 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_996
timestamp 1669390400
transform 1 0 112896 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1060
timestamp 1669390400
transform 1 0 120064 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1064
timestamp 1669390400
transform 1 0 120512 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1067
timestamp 1669390400
transform 1 0 120848 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1131
timestamp 1669390400
transform 1 0 128016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1135
timestamp 1669390400
transform 1 0 128464 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1138
timestamp 1669390400
transform 1 0 128800 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1202
timestamp 1669390400
transform 1 0 135968 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1206
timestamp 1669390400
transform 1 0 136416 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_1209
timestamp 1669390400
transform 1 0 136752 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1273
timestamp 1669390400
transform 1 0 143920 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1277
timestamp 1669390400
transform 1 0 144368 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_1280
timestamp 1669390400
transform 1 0 144704 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_1297
timestamp 1669390400
transform 1 0 146608 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_1301
timestamp 1669390400
transform 1 0 147056 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_1309
timestamp 1669390400
transform 1 0 147952 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1669390400
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1669390400
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1669390400
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1669390400
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1669390400
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1669390400
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1669390400
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1669390400
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_456
timestamp 1669390400
transform 1 0 52416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1669390400
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_463
timestamp 1669390400
transform 1 0 53200 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_527
timestamp 1669390400
transform 1 0 60368 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_531
timestamp 1669390400
transform 1 0 60816 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_534
timestamp 1669390400
transform 1 0 61152 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_598
timestamp 1669390400
transform 1 0 68320 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_602
timestamp 1669390400
transform 1 0 68768 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_605
timestamp 1669390400
transform 1 0 69104 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_669
timestamp 1669390400
transform 1 0 76272 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_673
timestamp 1669390400
transform 1 0 76720 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_676
timestamp 1669390400
transform 1 0 77056 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_740
timestamp 1669390400
transform 1 0 84224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_744
timestamp 1669390400
transform 1 0 84672 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_747
timestamp 1669390400
transform 1 0 85008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_811
timestamp 1669390400
transform 1 0 92176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_815
timestamp 1669390400
transform 1 0 92624 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_818
timestamp 1669390400
transform 1 0 92960 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_882
timestamp 1669390400
transform 1 0 100128 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_886
timestamp 1669390400
transform 1 0 100576 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_889
timestamp 1669390400
transform 1 0 100912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_896
timestamp 1669390400
transform 1 0 101696 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_928
timestamp 1669390400
transform 1 0 105280 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_944
timestamp 1669390400
transform 1 0 107072 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_952
timestamp 1669390400
transform 1 0 107968 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_956
timestamp 1669390400
transform 1 0 108416 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_960
timestamp 1669390400
transform 1 0 108864 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1024
timestamp 1669390400
transform 1 0 116032 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1028
timestamp 1669390400
transform 1 0 116480 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1031
timestamp 1669390400
transform 1 0 116816 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1095
timestamp 1669390400
transform 1 0 123984 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1099
timestamp 1669390400
transform 1 0 124432 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1102
timestamp 1669390400
transform 1 0 124768 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1166
timestamp 1669390400
transform 1 0 131936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1170
timestamp 1669390400
transform 1 0 132384 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_1173
timestamp 1669390400
transform 1 0 132720 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_1237
timestamp 1669390400
transform 1 0 139888 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1241
timestamp 1669390400
transform 1 0 140336 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_1244
timestamp 1669390400
transform 1 0 140672 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_1276
timestamp 1669390400
transform 1 0 144256 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_1279
timestamp 1669390400
transform 1 0 144592 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_1295
timestamp 1669390400
transform 1 0 146384 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_1311
timestamp 1669390400
transform 1 0 148176 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1669390400
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1669390400
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1669390400
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1669390400
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1669390400
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1669390400
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1669390400
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_421
timestamp 1669390400
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1669390400
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_428
timestamp 1669390400
transform 1 0 49280 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_492
timestamp 1669390400
transform 1 0 56448 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1669390400
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_499
timestamp 1669390400
transform 1 0 57232 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_563
timestamp 1669390400
transform 1 0 64400 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_567
timestamp 1669390400
transform 1 0 64848 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_570
timestamp 1669390400
transform 1 0 65184 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_634
timestamp 1669390400
transform 1 0 72352 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_638
timestamp 1669390400
transform 1 0 72800 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_641
timestamp 1669390400
transform 1 0 73136 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_705
timestamp 1669390400
transform 1 0 80304 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_709
timestamp 1669390400
transform 1 0 80752 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_712
timestamp 1669390400
transform 1 0 81088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_776
timestamp 1669390400
transform 1 0 88256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_780
timestamp 1669390400
transform 1 0 88704 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_783
timestamp 1669390400
transform 1 0 89040 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_847
timestamp 1669390400
transform 1 0 96208 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_851
timestamp 1669390400
transform 1 0 96656 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_854
timestamp 1669390400
transform 1 0 96992 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_870
timestamp 1669390400
transform 1 0 98784 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_878
timestamp 1669390400
transform 1 0 99680 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_880
timestamp 1669390400
transform 1 0 99904 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_887
timestamp 1669390400
transform 1 0 100688 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_919
timestamp 1669390400
transform 1 0 104272 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_925
timestamp 1669390400
transform 1 0 104944 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_989
timestamp 1669390400
transform 1 0 112112 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_993
timestamp 1669390400
transform 1 0 112560 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_996
timestamp 1669390400
transform 1 0 112896 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1060
timestamp 1669390400
transform 1 0 120064 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1064
timestamp 1669390400
transform 1 0 120512 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1067
timestamp 1669390400
transform 1 0 120848 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1131
timestamp 1669390400
transform 1 0 128016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1135
timestamp 1669390400
transform 1 0 128464 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1138
timestamp 1669390400
transform 1 0 128800 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_1202
timestamp 1669390400
transform 1 0 135968 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1206
timestamp 1669390400
transform 1 0 136416 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_1209
timestamp 1669390400
transform 1 0 136752 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_1273
timestamp 1669390400
transform 1 0 143920 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1277
timestamp 1669390400
transform 1 0 144368 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_1280
timestamp 1669390400
transform 1 0 144704 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_1295
timestamp 1669390400
transform 1 0 146384 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_1311
timestamp 1669390400
transform 1 0 148176 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1669390400
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1669390400
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1669390400
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1669390400
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1669390400
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1669390400
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1669390400
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1669390400
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1669390400
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1669390400
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_456
timestamp 1669390400
transform 1 0 52416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1669390400
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_463
timestamp 1669390400
transform 1 0 53200 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_527
timestamp 1669390400
transform 1 0 60368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_531
timestamp 1669390400
transform 1 0 60816 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_534
timestamp 1669390400
transform 1 0 61152 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_598
timestamp 1669390400
transform 1 0 68320 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_602
timestamp 1669390400
transform 1 0 68768 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_605
timestamp 1669390400
transform 1 0 69104 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_669
timestamp 1669390400
transform 1 0 76272 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_673
timestamp 1669390400
transform 1 0 76720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_676
timestamp 1669390400
transform 1 0 77056 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_740
timestamp 1669390400
transform 1 0 84224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_744
timestamp 1669390400
transform 1 0 84672 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_747
timestamp 1669390400
transform 1 0 85008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_811
timestamp 1669390400
transform 1 0 92176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_815
timestamp 1669390400
transform 1 0 92624 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_818
timestamp 1669390400
transform 1 0 92960 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_882
timestamp 1669390400
transform 1 0 100128 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_886
timestamp 1669390400
transform 1 0 100576 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_889
timestamp 1669390400
transform 1 0 100912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_896
timestamp 1669390400
transform 1 0 101696 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_928
timestamp 1669390400
transform 1 0 105280 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_944
timestamp 1669390400
transform 1 0 107072 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_952
timestamp 1669390400
transform 1 0 107968 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_956
timestamp 1669390400
transform 1 0 108416 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_960
timestamp 1669390400
transform 1 0 108864 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1024
timestamp 1669390400
transform 1 0 116032 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1028
timestamp 1669390400
transform 1 0 116480 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1031
timestamp 1669390400
transform 1 0 116816 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1095
timestamp 1669390400
transform 1 0 123984 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1099
timestamp 1669390400
transform 1 0 124432 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1102
timestamp 1669390400
transform 1 0 124768 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1166
timestamp 1669390400
transform 1 0 131936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1170
timestamp 1669390400
transform 1 0 132384 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_1173
timestamp 1669390400
transform 1 0 132720 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_1237
timestamp 1669390400
transform 1 0 139888 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1241
timestamp 1669390400
transform 1 0 140336 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_1244
timestamp 1669390400
transform 1 0 140672 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_1276
timestamp 1669390400
transform 1 0 144256 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_1279
timestamp 1669390400
transform 1 0 144592 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_1295
timestamp 1669390400
transform 1 0 146384 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_1311
timestamp 1669390400
transform 1 0 148176 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1669390400
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1669390400
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1669390400
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1669390400
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1669390400
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1669390400
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1669390400
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1669390400
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1669390400
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_421
timestamp 1669390400
transform 1 0 48496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1669390400
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_428
timestamp 1669390400
transform 1 0 49280 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_492
timestamp 1669390400
transform 1 0 56448 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_496
timestamp 1669390400
transform 1 0 56896 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_499
timestamp 1669390400
transform 1 0 57232 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_563
timestamp 1669390400
transform 1 0 64400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_567
timestamp 1669390400
transform 1 0 64848 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_570
timestamp 1669390400
transform 1 0 65184 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_634
timestamp 1669390400
transform 1 0 72352 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_638
timestamp 1669390400
transform 1 0 72800 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_641
timestamp 1669390400
transform 1 0 73136 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_705
timestamp 1669390400
transform 1 0 80304 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_709
timestamp 1669390400
transform 1 0 80752 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_712
timestamp 1669390400
transform 1 0 81088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_776
timestamp 1669390400
transform 1 0 88256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_780
timestamp 1669390400
transform 1 0 88704 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_783
timestamp 1669390400
transform 1 0 89040 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_847
timestamp 1669390400
transform 1 0 96208 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_851
timestamp 1669390400
transform 1 0 96656 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_854
timestamp 1669390400
transform 1 0 96992 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_918
timestamp 1669390400
transform 1 0 104160 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_922
timestamp 1669390400
transform 1 0 104608 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_925
timestamp 1669390400
transform 1 0 104944 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_989
timestamp 1669390400
transform 1 0 112112 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_993
timestamp 1669390400
transform 1 0 112560 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_996
timestamp 1669390400
transform 1 0 112896 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1060
timestamp 1669390400
transform 1 0 120064 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1064
timestamp 1669390400
transform 1 0 120512 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1067
timestamp 1669390400
transform 1 0 120848 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1131
timestamp 1669390400
transform 1 0 128016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1135
timestamp 1669390400
transform 1 0 128464 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1138
timestamp 1669390400
transform 1 0 128800 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1202
timestamp 1669390400
transform 1 0 135968 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1206
timestamp 1669390400
transform 1 0 136416 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_1209
timestamp 1669390400
transform 1 0 136752 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_1273
timestamp 1669390400
transform 1 0 143920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1277
timestamp 1669390400
transform 1 0 144368 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_1280
timestamp 1669390400
transform 1 0 144704 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_1312
timestamp 1669390400
transform 1 0 148288 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1669390400
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1669390400
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1669390400
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1669390400
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1669390400
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1669390400
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1669390400
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1669390400
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_456
timestamp 1669390400
transform 1 0 52416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_460
timestamp 1669390400
transform 1 0 52864 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_463
timestamp 1669390400
transform 1 0 53200 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_527
timestamp 1669390400
transform 1 0 60368 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_531
timestamp 1669390400
transform 1 0 60816 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_534
timestamp 1669390400
transform 1 0 61152 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_598
timestamp 1669390400
transform 1 0 68320 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_602
timestamp 1669390400
transform 1 0 68768 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_605
timestamp 1669390400
transform 1 0 69104 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_669
timestamp 1669390400
transform 1 0 76272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_673
timestamp 1669390400
transform 1 0 76720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_676
timestamp 1669390400
transform 1 0 77056 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_740
timestamp 1669390400
transform 1 0 84224 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_744
timestamp 1669390400
transform 1 0 84672 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_747
timestamp 1669390400
transform 1 0 85008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_811
timestamp 1669390400
transform 1 0 92176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_815
timestamp 1669390400
transform 1 0 92624 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_818
timestamp 1669390400
transform 1 0 92960 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_882
timestamp 1669390400
transform 1 0 100128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_886
timestamp 1669390400
transform 1 0 100576 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_889
timestamp 1669390400
transform 1 0 100912 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_953
timestamp 1669390400
transform 1 0 108080 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_957
timestamp 1669390400
transform 1 0 108528 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_960
timestamp 1669390400
transform 1 0 108864 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1024
timestamp 1669390400
transform 1 0 116032 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1028
timestamp 1669390400
transform 1 0 116480 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1031
timestamp 1669390400
transform 1 0 116816 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1095
timestamp 1669390400
transform 1 0 123984 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1099
timestamp 1669390400
transform 1 0 124432 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1102
timestamp 1669390400
transform 1 0 124768 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1166
timestamp 1669390400
transform 1 0 131936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1170
timestamp 1669390400
transform 1 0 132384 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_1173
timestamp 1669390400
transform 1 0 132720 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_1237
timestamp 1669390400
transform 1 0 139888 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1241
timestamp 1669390400
transform 1 0 140336 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_14_1244
timestamp 1669390400
transform 1 0 140672 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_1276
timestamp 1669390400
transform 1 0 144256 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_1279
timestamp 1669390400
transform 1 0 144592 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_1295
timestamp 1669390400
transform 1 0 146384 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_1311
timestamp 1669390400
transform 1 0 148176 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1669390400
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1669390400
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1669390400
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1669390400
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1669390400
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1669390400
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_421
timestamp 1669390400
transform 1 0 48496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1669390400
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_428
timestamp 1669390400
transform 1 0 49280 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_492
timestamp 1669390400
transform 1 0 56448 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1669390400
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_499
timestamp 1669390400
transform 1 0 57232 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_563
timestamp 1669390400
transform 1 0 64400 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_567
timestamp 1669390400
transform 1 0 64848 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_570
timestamp 1669390400
transform 1 0 65184 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_634
timestamp 1669390400
transform 1 0 72352 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_638
timestamp 1669390400
transform 1 0 72800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_641
timestamp 1669390400
transform 1 0 73136 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_705
timestamp 1669390400
transform 1 0 80304 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_709
timestamp 1669390400
transform 1 0 80752 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_712
timestamp 1669390400
transform 1 0 81088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_776
timestamp 1669390400
transform 1 0 88256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_780
timestamp 1669390400
transform 1 0 88704 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_783
timestamp 1669390400
transform 1 0 89040 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_847
timestamp 1669390400
transform 1 0 96208 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_851
timestamp 1669390400
transform 1 0 96656 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_854
timestamp 1669390400
transform 1 0 96992 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_918
timestamp 1669390400
transform 1 0 104160 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_922
timestamp 1669390400
transform 1 0 104608 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_925
timestamp 1669390400
transform 1 0 104944 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_989
timestamp 1669390400
transform 1 0 112112 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_993
timestamp 1669390400
transform 1 0 112560 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_996
timestamp 1669390400
transform 1 0 112896 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1060
timestamp 1669390400
transform 1 0 120064 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1064
timestamp 1669390400
transform 1 0 120512 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1067
timestamp 1669390400
transform 1 0 120848 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1131
timestamp 1669390400
transform 1 0 128016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1135
timestamp 1669390400
transform 1 0 128464 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1138
timestamp 1669390400
transform 1 0 128800 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_1202
timestamp 1669390400
transform 1 0 135968 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1206
timestamp 1669390400
transform 1 0 136416 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_1209
timestamp 1669390400
transform 1 0 136752 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_1273
timestamp 1669390400
transform 1 0 143920 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1277
timestamp 1669390400
transform 1 0 144368 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_1280
timestamp 1669390400
transform 1 0 144704 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_1295
timestamp 1669390400
transform 1 0 146384 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_1311
timestamp 1669390400
transform 1 0 148176 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1669390400
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1669390400
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1669390400
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1669390400
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1669390400
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1669390400
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_456
timestamp 1669390400
transform 1 0 52416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1669390400
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_463
timestamp 1669390400
transform 1 0 53200 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_527
timestamp 1669390400
transform 1 0 60368 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_531
timestamp 1669390400
transform 1 0 60816 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_534
timestamp 1669390400
transform 1 0 61152 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_598
timestamp 1669390400
transform 1 0 68320 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_602
timestamp 1669390400
transform 1 0 68768 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_605
timestamp 1669390400
transform 1 0 69104 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_669
timestamp 1669390400
transform 1 0 76272 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_673
timestamp 1669390400
transform 1 0 76720 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_676
timestamp 1669390400
transform 1 0 77056 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_740
timestamp 1669390400
transform 1 0 84224 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_744
timestamp 1669390400
transform 1 0 84672 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_747
timestamp 1669390400
transform 1 0 85008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_811
timestamp 1669390400
transform 1 0 92176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_815
timestamp 1669390400
transform 1 0 92624 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_818
timestamp 1669390400
transform 1 0 92960 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_882
timestamp 1669390400
transform 1 0 100128 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_886
timestamp 1669390400
transform 1 0 100576 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_889
timestamp 1669390400
transform 1 0 100912 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_953
timestamp 1669390400
transform 1 0 108080 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_957
timestamp 1669390400
transform 1 0 108528 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_960
timestamp 1669390400
transform 1 0 108864 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1024
timestamp 1669390400
transform 1 0 116032 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1028
timestamp 1669390400
transform 1 0 116480 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1031
timestamp 1669390400
transform 1 0 116816 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1095
timestamp 1669390400
transform 1 0 123984 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1099
timestamp 1669390400
transform 1 0 124432 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1102
timestamp 1669390400
transform 1 0 124768 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1166
timestamp 1669390400
transform 1 0 131936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1170
timestamp 1669390400
transform 1 0 132384 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_1173
timestamp 1669390400
transform 1 0 132720 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_1237
timestamp 1669390400
transform 1 0 139888 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1241
timestamp 1669390400
transform 1 0 140336 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_16_1244
timestamp 1669390400
transform 1 0 140672 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_1276
timestamp 1669390400
transform 1 0 144256 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1279
timestamp 1669390400
transform 1 0 144592 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_1295
timestamp 1669390400
transform 1 0 146384 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_1311
timestamp 1669390400
transform 1 0 148176 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1669390400
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1669390400
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1669390400
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1669390400
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1669390400
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1669390400
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1669390400
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_421
timestamp 1669390400
transform 1 0 48496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_425
timestamp 1669390400
transform 1 0 48944 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_428
timestamp 1669390400
transform 1 0 49280 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_492
timestamp 1669390400
transform 1 0 56448 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1669390400
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_499
timestamp 1669390400
transform 1 0 57232 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_563
timestamp 1669390400
transform 1 0 64400 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_567
timestamp 1669390400
transform 1 0 64848 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_570
timestamp 1669390400
transform 1 0 65184 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_634
timestamp 1669390400
transform 1 0 72352 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_638
timestamp 1669390400
transform 1 0 72800 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_641
timestamp 1669390400
transform 1 0 73136 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_705
timestamp 1669390400
transform 1 0 80304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_709
timestamp 1669390400
transform 1 0 80752 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_712
timestamp 1669390400
transform 1 0 81088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_776
timestamp 1669390400
transform 1 0 88256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_780
timestamp 1669390400
transform 1 0 88704 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_783
timestamp 1669390400
transform 1 0 89040 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_847
timestamp 1669390400
transform 1 0 96208 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_851
timestamp 1669390400
transform 1 0 96656 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_854
timestamp 1669390400
transform 1 0 96992 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_918
timestamp 1669390400
transform 1 0 104160 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_922
timestamp 1669390400
transform 1 0 104608 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_925
timestamp 1669390400
transform 1 0 104944 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_989
timestamp 1669390400
transform 1 0 112112 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_993
timestamp 1669390400
transform 1 0 112560 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_996
timestamp 1669390400
transform 1 0 112896 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1060
timestamp 1669390400
transform 1 0 120064 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1064
timestamp 1669390400
transform 1 0 120512 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1067
timestamp 1669390400
transform 1 0 120848 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1131
timestamp 1669390400
transform 1 0 128016 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1135
timestamp 1669390400
transform 1 0 128464 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1138
timestamp 1669390400
transform 1 0 128800 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_1202
timestamp 1669390400
transform 1 0 135968 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1206
timestamp 1669390400
transform 1 0 136416 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_1209
timestamp 1669390400
transform 1 0 136752 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_1273
timestamp 1669390400
transform 1 0 143920 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1277
timestamp 1669390400
transform 1 0 144368 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_1280
timestamp 1669390400
transform 1 0 144704 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_1295
timestamp 1669390400
transform 1 0 146384 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_1311
timestamp 1669390400
transform 1 0 148176 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1669390400
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1669390400
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1669390400
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1669390400
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1669390400
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1669390400
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1669390400
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_456
timestamp 1669390400
transform 1 0 52416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1669390400
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_463
timestamp 1669390400
transform 1 0 53200 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_527
timestamp 1669390400
transform 1 0 60368 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_531
timestamp 1669390400
transform 1 0 60816 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_534
timestamp 1669390400
transform 1 0 61152 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_598
timestamp 1669390400
transform 1 0 68320 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_602
timestamp 1669390400
transform 1 0 68768 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_605
timestamp 1669390400
transform 1 0 69104 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_669
timestamp 1669390400
transform 1 0 76272 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_673
timestamp 1669390400
transform 1 0 76720 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_676
timestamp 1669390400
transform 1 0 77056 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_740
timestamp 1669390400
transform 1 0 84224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_744
timestamp 1669390400
transform 1 0 84672 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_747
timestamp 1669390400
transform 1 0 85008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_811
timestamp 1669390400
transform 1 0 92176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_815
timestamp 1669390400
transform 1 0 92624 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_818
timestamp 1669390400
transform 1 0 92960 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_882
timestamp 1669390400
transform 1 0 100128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_886
timestamp 1669390400
transform 1 0 100576 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_889
timestamp 1669390400
transform 1 0 100912 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_953
timestamp 1669390400
transform 1 0 108080 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_957
timestamp 1669390400
transform 1 0 108528 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_960
timestamp 1669390400
transform 1 0 108864 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1024
timestamp 1669390400
transform 1 0 116032 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1028
timestamp 1669390400
transform 1 0 116480 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1031
timestamp 1669390400
transform 1 0 116816 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1095
timestamp 1669390400
transform 1 0 123984 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1099
timestamp 1669390400
transform 1 0 124432 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1102
timestamp 1669390400
transform 1 0 124768 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1166
timestamp 1669390400
transform 1 0 131936 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1170
timestamp 1669390400
transform 1 0 132384 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_1173
timestamp 1669390400
transform 1 0 132720 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_1237
timestamp 1669390400
transform 1 0 139888 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1241
timestamp 1669390400
transform 1 0 140336 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_18_1244
timestamp 1669390400
transform 1 0 140672 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_1276
timestamp 1669390400
transform 1 0 144256 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_1279
timestamp 1669390400
transform 1 0 144592 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_1295
timestamp 1669390400
transform 1 0 146384 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_1311
timestamp 1669390400
transform 1 0 148176 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1669390400
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1669390400
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1669390400
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1669390400
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1669390400
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1669390400
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1669390400
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_421
timestamp 1669390400
transform 1 0 48496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1669390400
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_428
timestamp 1669390400
transform 1 0 49280 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_492
timestamp 1669390400
transform 1 0 56448 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_496
timestamp 1669390400
transform 1 0 56896 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_499
timestamp 1669390400
transform 1 0 57232 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_563
timestamp 1669390400
transform 1 0 64400 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_567
timestamp 1669390400
transform 1 0 64848 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_570
timestamp 1669390400
transform 1 0 65184 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_634
timestamp 1669390400
transform 1 0 72352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_638
timestamp 1669390400
transform 1 0 72800 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_641
timestamp 1669390400
transform 1 0 73136 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_705
timestamp 1669390400
transform 1 0 80304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_709
timestamp 1669390400
transform 1 0 80752 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_712
timestamp 1669390400
transform 1 0 81088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_776
timestamp 1669390400
transform 1 0 88256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_780
timestamp 1669390400
transform 1 0 88704 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_783
timestamp 1669390400
transform 1 0 89040 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_847
timestamp 1669390400
transform 1 0 96208 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_851
timestamp 1669390400
transform 1 0 96656 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_854
timestamp 1669390400
transform 1 0 96992 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_918
timestamp 1669390400
transform 1 0 104160 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_922
timestamp 1669390400
transform 1 0 104608 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_925
timestamp 1669390400
transform 1 0 104944 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_957
timestamp 1669390400
transform 1 0 108528 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_973
timestamp 1669390400
transform 1 0 110320 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_975
timestamp 1669390400
transform 1 0 110544 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_978
timestamp 1669390400
transform 1 0 110880 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_986
timestamp 1669390400
transform 1 0 111776 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_996
timestamp 1669390400
transform 1 0 112896 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1060
timestamp 1669390400
transform 1 0 120064 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1064
timestamp 1669390400
transform 1 0 120512 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1067
timestamp 1669390400
transform 1 0 120848 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1131
timestamp 1669390400
transform 1 0 128016 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1135
timestamp 1669390400
transform 1 0 128464 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1138
timestamp 1669390400
transform 1 0 128800 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_1202
timestamp 1669390400
transform 1 0 135968 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1206
timestamp 1669390400
transform 1 0 136416 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_1209
timestamp 1669390400
transform 1 0 136752 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_1273
timestamp 1669390400
transform 1 0 143920 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1277
timestamp 1669390400
transform 1 0 144368 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_1280
timestamp 1669390400
transform 1 0 144704 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_1295
timestamp 1669390400
transform 1 0 146384 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_1311
timestamp 1669390400
transform 1 0 148176 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1669390400
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1669390400
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1669390400
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1669390400
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1669390400
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1669390400
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1669390400
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1669390400
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_456
timestamp 1669390400
transform 1 0 52416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_460
timestamp 1669390400
transform 1 0 52864 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_463
timestamp 1669390400
transform 1 0 53200 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_527
timestamp 1669390400
transform 1 0 60368 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_531
timestamp 1669390400
transform 1 0 60816 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_534
timestamp 1669390400
transform 1 0 61152 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_598
timestamp 1669390400
transform 1 0 68320 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_602
timestamp 1669390400
transform 1 0 68768 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_605
timestamp 1669390400
transform 1 0 69104 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_669
timestamp 1669390400
transform 1 0 76272 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_673
timestamp 1669390400
transform 1 0 76720 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_676
timestamp 1669390400
transform 1 0 77056 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_740
timestamp 1669390400
transform 1 0 84224 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_744
timestamp 1669390400
transform 1 0 84672 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_747
timestamp 1669390400
transform 1 0 85008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_811
timestamp 1669390400
transform 1 0 92176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_815
timestamp 1669390400
transform 1 0 92624 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_818
timestamp 1669390400
transform 1 0 92960 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_882
timestamp 1669390400
transform 1 0 100128 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_886
timestamp 1669390400
transform 1 0 100576 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_889
timestamp 1669390400
transform 1 0 100912 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_953
timestamp 1669390400
transform 1 0 108080 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_957
timestamp 1669390400
transform 1 0 108528 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_960
timestamp 1669390400
transform 1 0 108864 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1024
timestamp 1669390400
transform 1 0 116032 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1028
timestamp 1669390400
transform 1 0 116480 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1031
timestamp 1669390400
transform 1 0 116816 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1095
timestamp 1669390400
transform 1 0 123984 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1099
timestamp 1669390400
transform 1 0 124432 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1102
timestamp 1669390400
transform 1 0 124768 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1166
timestamp 1669390400
transform 1 0 131936 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1170
timestamp 1669390400
transform 1 0 132384 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_1173
timestamp 1669390400
transform 1 0 132720 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_1237
timestamp 1669390400
transform 1 0 139888 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1241
timestamp 1669390400
transform 1 0 140336 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_20_1244
timestamp 1669390400
transform 1 0 140672 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_1276
timestamp 1669390400
transform 1 0 144256 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_1279
timestamp 1669390400
transform 1 0 144592 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_1295
timestamp 1669390400
transform 1 0 146384 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_1311
timestamp 1669390400
transform 1 0 148176 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1669390400
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1669390400
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1669390400
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1669390400
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1669390400
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1669390400
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_421
timestamp 1669390400
transform 1 0 48496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1669390400
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_428
timestamp 1669390400
transform 1 0 49280 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_492
timestamp 1669390400
transform 1 0 56448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1669390400
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_499
timestamp 1669390400
transform 1 0 57232 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_563
timestamp 1669390400
transform 1 0 64400 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_567
timestamp 1669390400
transform 1 0 64848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_570
timestamp 1669390400
transform 1 0 65184 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_634
timestamp 1669390400
transform 1 0 72352 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_638
timestamp 1669390400
transform 1 0 72800 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_641
timestamp 1669390400
transform 1 0 73136 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_705
timestamp 1669390400
transform 1 0 80304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_709
timestamp 1669390400
transform 1 0 80752 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_712
timestamp 1669390400
transform 1 0 81088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_776
timestamp 1669390400
transform 1 0 88256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_780
timestamp 1669390400
transform 1 0 88704 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_783
timestamp 1669390400
transform 1 0 89040 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_847
timestamp 1669390400
transform 1 0 96208 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_851
timestamp 1669390400
transform 1 0 96656 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_854
timestamp 1669390400
transform 1 0 96992 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_918
timestamp 1669390400
transform 1 0 104160 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_922
timestamp 1669390400
transform 1 0 104608 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_925
timestamp 1669390400
transform 1 0 104944 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_989
timestamp 1669390400
transform 1 0 112112 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_993
timestamp 1669390400
transform 1 0 112560 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_996
timestamp 1669390400
transform 1 0 112896 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1060
timestamp 1669390400
transform 1 0 120064 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1064
timestamp 1669390400
transform 1 0 120512 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1067
timestamp 1669390400
transform 1 0 120848 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1131
timestamp 1669390400
transform 1 0 128016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1135
timestamp 1669390400
transform 1 0 128464 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1138
timestamp 1669390400
transform 1 0 128800 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1202
timestamp 1669390400
transform 1 0 135968 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1206
timestamp 1669390400
transform 1 0 136416 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_1209
timestamp 1669390400
transform 1 0 136752 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_1273
timestamp 1669390400
transform 1 0 143920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1277
timestamp 1669390400
transform 1 0 144368 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_1280
timestamp 1669390400
transform 1 0 144704 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_1312
timestamp 1669390400
transform 1 0 148288 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1669390400
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1669390400
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1669390400
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1669390400
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1669390400
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1669390400
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1669390400
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1669390400
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1669390400
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1669390400
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_456
timestamp 1669390400
transform 1 0 52416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_460
timestamp 1669390400
transform 1 0 52864 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_463
timestamp 1669390400
transform 1 0 53200 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_527
timestamp 1669390400
transform 1 0 60368 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_531
timestamp 1669390400
transform 1 0 60816 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_534
timestamp 1669390400
transform 1 0 61152 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_598
timestamp 1669390400
transform 1 0 68320 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_602
timestamp 1669390400
transform 1 0 68768 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_605
timestamp 1669390400
transform 1 0 69104 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_669
timestamp 1669390400
transform 1 0 76272 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_673
timestamp 1669390400
transform 1 0 76720 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_676
timestamp 1669390400
transform 1 0 77056 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_740
timestamp 1669390400
transform 1 0 84224 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_744
timestamp 1669390400
transform 1 0 84672 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_747
timestamp 1669390400
transform 1 0 85008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_811
timestamp 1669390400
transform 1 0 92176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_815
timestamp 1669390400
transform 1 0 92624 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_818
timestamp 1669390400
transform 1 0 92960 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_882
timestamp 1669390400
transform 1 0 100128 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_886
timestamp 1669390400
transform 1 0 100576 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_889
timestamp 1669390400
transform 1 0 100912 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_953
timestamp 1669390400
transform 1 0 108080 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_957
timestamp 1669390400
transform 1 0 108528 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_960
timestamp 1669390400
transform 1 0 108864 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1024
timestamp 1669390400
transform 1 0 116032 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1028
timestamp 1669390400
transform 1 0 116480 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1031
timestamp 1669390400
transform 1 0 116816 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1095
timestamp 1669390400
transform 1 0 123984 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1099
timestamp 1669390400
transform 1 0 124432 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1102
timestamp 1669390400
transform 1 0 124768 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1166
timestamp 1669390400
transform 1 0 131936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1170
timestamp 1669390400
transform 1 0 132384 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_1173
timestamp 1669390400
transform 1 0 132720 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_1237
timestamp 1669390400
transform 1 0 139888 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1241
timestamp 1669390400
transform 1 0 140336 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_1244
timestamp 1669390400
transform 1 0 140672 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_1276
timestamp 1669390400
transform 1 0 144256 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_1279
timestamp 1669390400
transform 1 0 144592 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_1295
timestamp 1669390400
transform 1 0 146384 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_1311
timestamp 1669390400
transform 1 0 148176 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_66
timestamp 1669390400
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1669390400
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1669390400
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1669390400
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1669390400
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1669390400
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_421
timestamp 1669390400
transform 1 0 48496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_425
timestamp 1669390400
transform 1 0 48944 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_428
timestamp 1669390400
transform 1 0 49280 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_492
timestamp 1669390400
transform 1 0 56448 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1669390400
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_499
timestamp 1669390400
transform 1 0 57232 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_563
timestamp 1669390400
transform 1 0 64400 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_567
timestamp 1669390400
transform 1 0 64848 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_570
timestamp 1669390400
transform 1 0 65184 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_634
timestamp 1669390400
transform 1 0 72352 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_638
timestamp 1669390400
transform 1 0 72800 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_641
timestamp 1669390400
transform 1 0 73136 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_705
timestamp 1669390400
transform 1 0 80304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_709
timestamp 1669390400
transform 1 0 80752 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_712
timestamp 1669390400
transform 1 0 81088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_776
timestamp 1669390400
transform 1 0 88256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_780
timestamp 1669390400
transform 1 0 88704 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_783
timestamp 1669390400
transform 1 0 89040 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_847
timestamp 1669390400
transform 1 0 96208 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_851
timestamp 1669390400
transform 1 0 96656 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_854
timestamp 1669390400
transform 1 0 96992 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_918
timestamp 1669390400
transform 1 0 104160 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_922
timestamp 1669390400
transform 1 0 104608 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_925
timestamp 1669390400
transform 1 0 104944 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_989
timestamp 1669390400
transform 1 0 112112 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_993
timestamp 1669390400
transform 1 0 112560 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_996
timestamp 1669390400
transform 1 0 112896 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1060
timestamp 1669390400
transform 1 0 120064 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1064
timestamp 1669390400
transform 1 0 120512 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1067
timestamp 1669390400
transform 1 0 120848 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1131
timestamp 1669390400
transform 1 0 128016 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1135
timestamp 1669390400
transform 1 0 128464 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1138
timestamp 1669390400
transform 1 0 128800 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_1202
timestamp 1669390400
transform 1 0 135968 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1206
timestamp 1669390400
transform 1 0 136416 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_1209
timestamp 1669390400
transform 1 0 136752 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_1273
timestamp 1669390400
transform 1 0 143920 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1277
timestamp 1669390400
transform 1 0 144368 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_1280
timestamp 1669390400
transform 1 0 144704 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_1295
timestamp 1669390400
transform 1 0 146384 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_1311
timestamp 1669390400
transform 1 0 148176 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1669390400
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1669390400
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1669390400
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1669390400
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1669390400
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1669390400
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1669390400
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_456
timestamp 1669390400
transform 1 0 52416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_460
timestamp 1669390400
transform 1 0 52864 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_463
timestamp 1669390400
transform 1 0 53200 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_527
timestamp 1669390400
transform 1 0 60368 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_531
timestamp 1669390400
transform 1 0 60816 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_534
timestamp 1669390400
transform 1 0 61152 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_598
timestamp 1669390400
transform 1 0 68320 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_602
timestamp 1669390400
transform 1 0 68768 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_605
timestamp 1669390400
transform 1 0 69104 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_669
timestamp 1669390400
transform 1 0 76272 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_673
timestamp 1669390400
transform 1 0 76720 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_676
timestamp 1669390400
transform 1 0 77056 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_740
timestamp 1669390400
transform 1 0 84224 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_744
timestamp 1669390400
transform 1 0 84672 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_747
timestamp 1669390400
transform 1 0 85008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_811
timestamp 1669390400
transform 1 0 92176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_815
timestamp 1669390400
transform 1 0 92624 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_818
timestamp 1669390400
transform 1 0 92960 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_882
timestamp 1669390400
transform 1 0 100128 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_886
timestamp 1669390400
transform 1 0 100576 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_889
timestamp 1669390400
transform 1 0 100912 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_953
timestamp 1669390400
transform 1 0 108080 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_957
timestamp 1669390400
transform 1 0 108528 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_960
timestamp 1669390400
transform 1 0 108864 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1024
timestamp 1669390400
transform 1 0 116032 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1028
timestamp 1669390400
transform 1 0 116480 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1031
timestamp 1669390400
transform 1 0 116816 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1095
timestamp 1669390400
transform 1 0 123984 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1099
timestamp 1669390400
transform 1 0 124432 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1102
timestamp 1669390400
transform 1 0 124768 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1166
timestamp 1669390400
transform 1 0 131936 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1170
timestamp 1669390400
transform 1 0 132384 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_1173
timestamp 1669390400
transform 1 0 132720 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_1237
timestamp 1669390400
transform 1 0 139888 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1241
timestamp 1669390400
transform 1 0 140336 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_1244
timestamp 1669390400
transform 1 0 140672 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_1276
timestamp 1669390400
transform 1 0 144256 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_1279
timestamp 1669390400
transform 1 0 144592 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_1295
timestamp 1669390400
transform 1 0 146384 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_1311
timestamp 1669390400
transform 1 0 148176 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_66
timestamp 1669390400
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1669390400
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1669390400
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1669390400
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1669390400
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1669390400
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_421
timestamp 1669390400
transform 1 0 48496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_425
timestamp 1669390400
transform 1 0 48944 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_428
timestamp 1669390400
transform 1 0 49280 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_492
timestamp 1669390400
transform 1 0 56448 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1669390400
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_499
timestamp 1669390400
transform 1 0 57232 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_563
timestamp 1669390400
transform 1 0 64400 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_567
timestamp 1669390400
transform 1 0 64848 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_570
timestamp 1669390400
transform 1 0 65184 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_634
timestamp 1669390400
transform 1 0 72352 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_638
timestamp 1669390400
transform 1 0 72800 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_641
timestamp 1669390400
transform 1 0 73136 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_705
timestamp 1669390400
transform 1 0 80304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_709
timestamp 1669390400
transform 1 0 80752 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_712
timestamp 1669390400
transform 1 0 81088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_776
timestamp 1669390400
transform 1 0 88256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_780
timestamp 1669390400
transform 1 0 88704 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_783
timestamp 1669390400
transform 1 0 89040 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_847
timestamp 1669390400
transform 1 0 96208 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_851
timestamp 1669390400
transform 1 0 96656 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_854
timestamp 1669390400
transform 1 0 96992 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_918
timestamp 1669390400
transform 1 0 104160 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_922
timestamp 1669390400
transform 1 0 104608 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_925
timestamp 1669390400
transform 1 0 104944 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_989
timestamp 1669390400
transform 1 0 112112 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_993
timestamp 1669390400
transform 1 0 112560 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_996
timestamp 1669390400
transform 1 0 112896 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1060
timestamp 1669390400
transform 1 0 120064 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1064
timestamp 1669390400
transform 1 0 120512 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1067
timestamp 1669390400
transform 1 0 120848 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1131
timestamp 1669390400
transform 1 0 128016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1135
timestamp 1669390400
transform 1 0 128464 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1138
timestamp 1669390400
transform 1 0 128800 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_1202
timestamp 1669390400
transform 1 0 135968 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1206
timestamp 1669390400
transform 1 0 136416 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_1209
timestamp 1669390400
transform 1 0 136752 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_1273
timestamp 1669390400
transform 1 0 143920 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1277
timestamp 1669390400
transform 1 0 144368 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_1280
timestamp 1669390400
transform 1 0 144704 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_1295
timestamp 1669390400
transform 1 0 146384 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_1311
timestamp 1669390400
transform 1 0 148176 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1669390400
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1669390400
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1669390400
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1669390400
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1669390400
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1669390400
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1669390400
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1669390400
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_456
timestamp 1669390400
transform 1 0 52416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_460
timestamp 1669390400
transform 1 0 52864 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_463
timestamp 1669390400
transform 1 0 53200 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_527
timestamp 1669390400
transform 1 0 60368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_531
timestamp 1669390400
transform 1 0 60816 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_534
timestamp 1669390400
transform 1 0 61152 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_598
timestamp 1669390400
transform 1 0 68320 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_602
timestamp 1669390400
transform 1 0 68768 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_605
timestamp 1669390400
transform 1 0 69104 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_669
timestamp 1669390400
transform 1 0 76272 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_673
timestamp 1669390400
transform 1 0 76720 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_676
timestamp 1669390400
transform 1 0 77056 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_740
timestamp 1669390400
transform 1 0 84224 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_744
timestamp 1669390400
transform 1 0 84672 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_747
timestamp 1669390400
transform 1 0 85008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_811
timestamp 1669390400
transform 1 0 92176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_815
timestamp 1669390400
transform 1 0 92624 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_818
timestamp 1669390400
transform 1 0 92960 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_882
timestamp 1669390400
transform 1 0 100128 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_886
timestamp 1669390400
transform 1 0 100576 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_889
timestamp 1669390400
transform 1 0 100912 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_953
timestamp 1669390400
transform 1 0 108080 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_957
timestamp 1669390400
transform 1 0 108528 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_960
timestamp 1669390400
transform 1 0 108864 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1024
timestamp 1669390400
transform 1 0 116032 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1028
timestamp 1669390400
transform 1 0 116480 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1031
timestamp 1669390400
transform 1 0 116816 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1095
timestamp 1669390400
transform 1 0 123984 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1099
timestamp 1669390400
transform 1 0 124432 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1102
timestamp 1669390400
transform 1 0 124768 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1166
timestamp 1669390400
transform 1 0 131936 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1170
timestamp 1669390400
transform 1 0 132384 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_1173
timestamp 1669390400
transform 1 0 132720 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_1237
timestamp 1669390400
transform 1 0 139888 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1241
timestamp 1669390400
transform 1 0 140336 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_1244
timestamp 1669390400
transform 1 0 140672 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_1276
timestamp 1669390400
transform 1 0 144256 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_1279
timestamp 1669390400
transform 1 0 144592 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_1295
timestamp 1669390400
transform 1 0 146384 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_1311
timestamp 1669390400
transform 1 0 148176 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_66
timestamp 1669390400
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1669390400
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1669390400
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1669390400
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1669390400
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1669390400
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_421
timestamp 1669390400
transform 1 0 48496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_425
timestamp 1669390400
transform 1 0 48944 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_428
timestamp 1669390400
transform 1 0 49280 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_492
timestamp 1669390400
transform 1 0 56448 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_496
timestamp 1669390400
transform 1 0 56896 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_499
timestamp 1669390400
transform 1 0 57232 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_563
timestamp 1669390400
transform 1 0 64400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_567
timestamp 1669390400
transform 1 0 64848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_570
timestamp 1669390400
transform 1 0 65184 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_634
timestamp 1669390400
transform 1 0 72352 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_638
timestamp 1669390400
transform 1 0 72800 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_641
timestamp 1669390400
transform 1 0 73136 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_705
timestamp 1669390400
transform 1 0 80304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_709
timestamp 1669390400
transform 1 0 80752 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_712
timestamp 1669390400
transform 1 0 81088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_776
timestamp 1669390400
transform 1 0 88256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_780
timestamp 1669390400
transform 1 0 88704 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_783
timestamp 1669390400
transform 1 0 89040 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_847
timestamp 1669390400
transform 1 0 96208 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_851
timestamp 1669390400
transform 1 0 96656 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_854
timestamp 1669390400
transform 1 0 96992 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_918
timestamp 1669390400
transform 1 0 104160 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_922
timestamp 1669390400
transform 1 0 104608 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_925
timestamp 1669390400
transform 1 0 104944 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_989
timestamp 1669390400
transform 1 0 112112 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_993
timestamp 1669390400
transform 1 0 112560 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_996
timestamp 1669390400
transform 1 0 112896 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1060
timestamp 1669390400
transform 1 0 120064 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1064
timestamp 1669390400
transform 1 0 120512 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1067
timestamp 1669390400
transform 1 0 120848 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1131
timestamp 1669390400
transform 1 0 128016 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1135
timestamp 1669390400
transform 1 0 128464 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1138
timestamp 1669390400
transform 1 0 128800 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_1202
timestamp 1669390400
transform 1 0 135968 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1206
timestamp 1669390400
transform 1 0 136416 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_1209
timestamp 1669390400
transform 1 0 136752 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_1273
timestamp 1669390400
transform 1 0 143920 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1277
timestamp 1669390400
transform 1 0 144368 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_1280
timestamp 1669390400
transform 1 0 144704 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_1295
timestamp 1669390400
transform 1 0 146384 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_1311
timestamp 1669390400
transform 1 0 148176 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1669390400
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1669390400
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1669390400
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1669390400
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1669390400
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1669390400
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1669390400
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1669390400
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_456
timestamp 1669390400
transform 1 0 52416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_460
timestamp 1669390400
transform 1 0 52864 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_463
timestamp 1669390400
transform 1 0 53200 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_527
timestamp 1669390400
transform 1 0 60368 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_531
timestamp 1669390400
transform 1 0 60816 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_534
timestamp 1669390400
transform 1 0 61152 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_598
timestamp 1669390400
transform 1 0 68320 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_602
timestamp 1669390400
transform 1 0 68768 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_605
timestamp 1669390400
transform 1 0 69104 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_669
timestamp 1669390400
transform 1 0 76272 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_673
timestamp 1669390400
transform 1 0 76720 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_676
timestamp 1669390400
transform 1 0 77056 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_740
timestamp 1669390400
transform 1 0 84224 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_744
timestamp 1669390400
transform 1 0 84672 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_747
timestamp 1669390400
transform 1 0 85008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_811
timestamp 1669390400
transform 1 0 92176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_815
timestamp 1669390400
transform 1 0 92624 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_818
timestamp 1669390400
transform 1 0 92960 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_882
timestamp 1669390400
transform 1 0 100128 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_886
timestamp 1669390400
transform 1 0 100576 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_889
timestamp 1669390400
transform 1 0 100912 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_953
timestamp 1669390400
transform 1 0 108080 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_957
timestamp 1669390400
transform 1 0 108528 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_960
timestamp 1669390400
transform 1 0 108864 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1024
timestamp 1669390400
transform 1 0 116032 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1028
timestamp 1669390400
transform 1 0 116480 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1031
timestamp 1669390400
transform 1 0 116816 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1095
timestamp 1669390400
transform 1 0 123984 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1099
timestamp 1669390400
transform 1 0 124432 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1102
timestamp 1669390400
transform 1 0 124768 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1166
timestamp 1669390400
transform 1 0 131936 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1170
timestamp 1669390400
transform 1 0 132384 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_1173
timestamp 1669390400
transform 1 0 132720 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_1237
timestamp 1669390400
transform 1 0 139888 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1241
timestamp 1669390400
transform 1 0 140336 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_1244
timestamp 1669390400
transform 1 0 140672 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_1276
timestamp 1669390400
transform 1 0 144256 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_1279
timestamp 1669390400
transform 1 0 144592 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_1295
timestamp 1669390400
transform 1 0 146384 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_1311
timestamp 1669390400
transform 1 0 148176 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1669390400
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1669390400
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1669390400
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1669390400
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1669390400
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_421
timestamp 1669390400
transform 1 0 48496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1669390400
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_428
timestamp 1669390400
transform 1 0 49280 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_492
timestamp 1669390400
transform 1 0 56448 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_496
timestamp 1669390400
transform 1 0 56896 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_499
timestamp 1669390400
transform 1 0 57232 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_563
timestamp 1669390400
transform 1 0 64400 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_567
timestamp 1669390400
transform 1 0 64848 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_570
timestamp 1669390400
transform 1 0 65184 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_634
timestamp 1669390400
transform 1 0 72352 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_638
timestamp 1669390400
transform 1 0 72800 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_641
timestamp 1669390400
transform 1 0 73136 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_705
timestamp 1669390400
transform 1 0 80304 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_709
timestamp 1669390400
transform 1 0 80752 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_712
timestamp 1669390400
transform 1 0 81088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_776
timestamp 1669390400
transform 1 0 88256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_780
timestamp 1669390400
transform 1 0 88704 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_783
timestamp 1669390400
transform 1 0 89040 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_847
timestamp 1669390400
transform 1 0 96208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_851
timestamp 1669390400
transform 1 0 96656 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_854
timestamp 1669390400
transform 1 0 96992 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_918
timestamp 1669390400
transform 1 0 104160 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_922
timestamp 1669390400
transform 1 0 104608 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_925
timestamp 1669390400
transform 1 0 104944 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_989
timestamp 1669390400
transform 1 0 112112 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_993
timestamp 1669390400
transform 1 0 112560 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_996
timestamp 1669390400
transform 1 0 112896 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1060
timestamp 1669390400
transform 1 0 120064 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1064
timestamp 1669390400
transform 1 0 120512 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1067
timestamp 1669390400
transform 1 0 120848 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1131
timestamp 1669390400
transform 1 0 128016 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1135
timestamp 1669390400
transform 1 0 128464 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1138
timestamp 1669390400
transform 1 0 128800 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1202
timestamp 1669390400
transform 1 0 135968 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1206
timestamp 1669390400
transform 1 0 136416 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_1209
timestamp 1669390400
transform 1 0 136752 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_1273
timestamp 1669390400
transform 1 0 143920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1277
timestamp 1669390400
transform 1 0 144368 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_1280
timestamp 1669390400
transform 1 0 144704 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_1312
timestamp 1669390400
transform 1 0 148288 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1669390400
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1669390400
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1669390400
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1669390400
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1669390400
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1669390400
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1669390400
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_456
timestamp 1669390400
transform 1 0 52416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_460
timestamp 1669390400
transform 1 0 52864 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_463
timestamp 1669390400
transform 1 0 53200 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_527
timestamp 1669390400
transform 1 0 60368 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_531
timestamp 1669390400
transform 1 0 60816 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_534
timestamp 1669390400
transform 1 0 61152 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_598
timestamp 1669390400
transform 1 0 68320 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_602
timestamp 1669390400
transform 1 0 68768 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_605
timestamp 1669390400
transform 1 0 69104 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_669
timestamp 1669390400
transform 1 0 76272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_673
timestamp 1669390400
transform 1 0 76720 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_676
timestamp 1669390400
transform 1 0 77056 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_740
timestamp 1669390400
transform 1 0 84224 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_744
timestamp 1669390400
transform 1 0 84672 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_747
timestamp 1669390400
transform 1 0 85008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_811
timestamp 1669390400
transform 1 0 92176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_815
timestamp 1669390400
transform 1 0 92624 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_818
timestamp 1669390400
transform 1 0 92960 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_882
timestamp 1669390400
transform 1 0 100128 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_886
timestamp 1669390400
transform 1 0 100576 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_889
timestamp 1669390400
transform 1 0 100912 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_953
timestamp 1669390400
transform 1 0 108080 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_957
timestamp 1669390400
transform 1 0 108528 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_960
timestamp 1669390400
transform 1 0 108864 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1024
timestamp 1669390400
transform 1 0 116032 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1028
timestamp 1669390400
transform 1 0 116480 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1031
timestamp 1669390400
transform 1 0 116816 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1095
timestamp 1669390400
transform 1 0 123984 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1099
timestamp 1669390400
transform 1 0 124432 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1102
timestamp 1669390400
transform 1 0 124768 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1166
timestamp 1669390400
transform 1 0 131936 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1170
timestamp 1669390400
transform 1 0 132384 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_1173
timestamp 1669390400
transform 1 0 132720 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_1237
timestamp 1669390400
transform 1 0 139888 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1241
timestamp 1669390400
transform 1 0 140336 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_30_1244
timestamp 1669390400
transform 1 0 140672 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_1276
timestamp 1669390400
transform 1 0 144256 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_1279
timestamp 1669390400
transform 1 0 144592 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_1295
timestamp 1669390400
transform 1 0 146384 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_1311
timestamp 1669390400
transform 1 0 148176 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1669390400
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1669390400
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1669390400
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1669390400
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1669390400
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1669390400
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1669390400
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1669390400
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1669390400
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1669390400
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_421
timestamp 1669390400
transform 1 0 48496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1669390400
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_428
timestamp 1669390400
transform 1 0 49280 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_492
timestamp 1669390400
transform 1 0 56448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1669390400
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_499
timestamp 1669390400
transform 1 0 57232 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_563
timestamp 1669390400
transform 1 0 64400 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_567
timestamp 1669390400
transform 1 0 64848 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_570
timestamp 1669390400
transform 1 0 65184 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_634
timestamp 1669390400
transform 1 0 72352 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_638
timestamp 1669390400
transform 1 0 72800 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_641
timestamp 1669390400
transform 1 0 73136 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_705
timestamp 1669390400
transform 1 0 80304 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_709
timestamp 1669390400
transform 1 0 80752 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_712
timestamp 1669390400
transform 1 0 81088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_776
timestamp 1669390400
transform 1 0 88256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_780
timestamp 1669390400
transform 1 0 88704 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_783
timestamp 1669390400
transform 1 0 89040 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_847
timestamp 1669390400
transform 1 0 96208 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_851
timestamp 1669390400
transform 1 0 96656 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_854
timestamp 1669390400
transform 1 0 96992 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_918
timestamp 1669390400
transform 1 0 104160 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_922
timestamp 1669390400
transform 1 0 104608 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_925
timestamp 1669390400
transform 1 0 104944 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_989
timestamp 1669390400
transform 1 0 112112 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_993
timestamp 1669390400
transform 1 0 112560 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_996
timestamp 1669390400
transform 1 0 112896 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1060
timestamp 1669390400
transform 1 0 120064 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1064
timestamp 1669390400
transform 1 0 120512 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1067
timestamp 1669390400
transform 1 0 120848 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1131
timestamp 1669390400
transform 1 0 128016 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1135
timestamp 1669390400
transform 1 0 128464 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1138
timestamp 1669390400
transform 1 0 128800 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_1202
timestamp 1669390400
transform 1 0 135968 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1206
timestamp 1669390400
transform 1 0 136416 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_1209
timestamp 1669390400
transform 1 0 136752 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_1273
timestamp 1669390400
transform 1 0 143920 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1277
timestamp 1669390400
transform 1 0 144368 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_1280
timestamp 1669390400
transform 1 0 144704 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_1295
timestamp 1669390400
transform 1 0 146384 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_1311
timestamp 1669390400
transform 1 0 148176 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1669390400
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1669390400
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1669390400
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_243
timestamp 1669390400
transform 1 0 28560 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_247
timestamp 1669390400
transform 1 0 29008 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1669390400
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1669390400
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1669390400
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1669390400
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_456
timestamp 1669390400
transform 1 0 52416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1669390400
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_463
timestamp 1669390400
transform 1 0 53200 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_527
timestamp 1669390400
transform 1 0 60368 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_531
timestamp 1669390400
transform 1 0 60816 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_534
timestamp 1669390400
transform 1 0 61152 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_598
timestamp 1669390400
transform 1 0 68320 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_602
timestamp 1669390400
transform 1 0 68768 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_605
timestamp 1669390400
transform 1 0 69104 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_669
timestamp 1669390400
transform 1 0 76272 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_673
timestamp 1669390400
transform 1 0 76720 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_676
timestamp 1669390400
transform 1 0 77056 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_740
timestamp 1669390400
transform 1 0 84224 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_744
timestamp 1669390400
transform 1 0 84672 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_747
timestamp 1669390400
transform 1 0 85008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_811
timestamp 1669390400
transform 1 0 92176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_815
timestamp 1669390400
transform 1 0 92624 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_818
timestamp 1669390400
transform 1 0 92960 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_882
timestamp 1669390400
transform 1 0 100128 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_886
timestamp 1669390400
transform 1 0 100576 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_889
timestamp 1669390400
transform 1 0 100912 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_953
timestamp 1669390400
transform 1 0 108080 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_957
timestamp 1669390400
transform 1 0 108528 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_960
timestamp 1669390400
transform 1 0 108864 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1024
timestamp 1669390400
transform 1 0 116032 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1028
timestamp 1669390400
transform 1 0 116480 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1031
timestamp 1669390400
transform 1 0 116816 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1095
timestamp 1669390400
transform 1 0 123984 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1099
timestamp 1669390400
transform 1 0 124432 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1102
timestamp 1669390400
transform 1 0 124768 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1166
timestamp 1669390400
transform 1 0 131936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1170
timestamp 1669390400
transform 1 0 132384 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_1173
timestamp 1669390400
transform 1 0 132720 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_1237
timestamp 1669390400
transform 1 0 139888 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1241
timestamp 1669390400
transform 1 0 140336 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_1244
timestamp 1669390400
transform 1 0 140672 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_1276
timestamp 1669390400
transform 1 0 144256 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_1279
timestamp 1669390400
transform 1 0 144592 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_1295
timestamp 1669390400
transform 1 0 146384 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_1311
timestamp 1669390400
transform 1 0 148176 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1669390400
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1669390400
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1669390400
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1669390400
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_208
timestamp 1669390400
transform 1 0 24640 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1669390400
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1669390400
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1669390400
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_421
timestamp 1669390400
transform 1 0 48496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1669390400
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_428
timestamp 1669390400
transform 1 0 49280 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_492
timestamp 1669390400
transform 1 0 56448 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1669390400
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_499
timestamp 1669390400
transform 1 0 57232 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_563
timestamp 1669390400
transform 1 0 64400 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_567
timestamp 1669390400
transform 1 0 64848 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_570
timestamp 1669390400
transform 1 0 65184 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_634
timestamp 1669390400
transform 1 0 72352 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_638
timestamp 1669390400
transform 1 0 72800 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_641
timestamp 1669390400
transform 1 0 73136 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_705
timestamp 1669390400
transform 1 0 80304 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_709
timestamp 1669390400
transform 1 0 80752 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_712
timestamp 1669390400
transform 1 0 81088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_776
timestamp 1669390400
transform 1 0 88256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_780
timestamp 1669390400
transform 1 0 88704 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_783
timestamp 1669390400
transform 1 0 89040 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_847
timestamp 1669390400
transform 1 0 96208 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_851
timestamp 1669390400
transform 1 0 96656 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_854
timestamp 1669390400
transform 1 0 96992 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_918
timestamp 1669390400
transform 1 0 104160 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_922
timestamp 1669390400
transform 1 0 104608 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_925
timestamp 1669390400
transform 1 0 104944 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_989
timestamp 1669390400
transform 1 0 112112 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_993
timestamp 1669390400
transform 1 0 112560 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_996
timestamp 1669390400
transform 1 0 112896 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1060
timestamp 1669390400
transform 1 0 120064 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1064
timestamp 1669390400
transform 1 0 120512 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1067
timestamp 1669390400
transform 1 0 120848 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1131
timestamp 1669390400
transform 1 0 128016 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1135
timestamp 1669390400
transform 1 0 128464 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1138
timestamp 1669390400
transform 1 0 128800 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_1202
timestamp 1669390400
transform 1 0 135968 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1206
timestamp 1669390400
transform 1 0 136416 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_1209
timestamp 1669390400
transform 1 0 136752 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_1273
timestamp 1669390400
transform 1 0 143920 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1277
timestamp 1669390400
transform 1 0 144368 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_1280
timestamp 1669390400
transform 1 0 144704 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_1295
timestamp 1669390400
transform 1 0 146384 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_1311
timestamp 1669390400
transform 1 0 148176 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1669390400
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1669390400
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_172
timestamp 1669390400
transform 1 0 20608 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_243
timestamp 1669390400
transform 1 0 28560 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1669390400
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1669390400
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1669390400
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_456
timestamp 1669390400
transform 1 0 52416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1669390400
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_463
timestamp 1669390400
transform 1 0 53200 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_527
timestamp 1669390400
transform 1 0 60368 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_531
timestamp 1669390400
transform 1 0 60816 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_534
timestamp 1669390400
transform 1 0 61152 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_598
timestamp 1669390400
transform 1 0 68320 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_602
timestamp 1669390400
transform 1 0 68768 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_605
timestamp 1669390400
transform 1 0 69104 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_669
timestamp 1669390400
transform 1 0 76272 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_673
timestamp 1669390400
transform 1 0 76720 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_676
timestamp 1669390400
transform 1 0 77056 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_740
timestamp 1669390400
transform 1 0 84224 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_744
timestamp 1669390400
transform 1 0 84672 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_747
timestamp 1669390400
transform 1 0 85008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_811
timestamp 1669390400
transform 1 0 92176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_815
timestamp 1669390400
transform 1 0 92624 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_818
timestamp 1669390400
transform 1 0 92960 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_882
timestamp 1669390400
transform 1 0 100128 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_886
timestamp 1669390400
transform 1 0 100576 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_889
timestamp 1669390400
transform 1 0 100912 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_953
timestamp 1669390400
transform 1 0 108080 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_957
timestamp 1669390400
transform 1 0 108528 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_960
timestamp 1669390400
transform 1 0 108864 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1024
timestamp 1669390400
transform 1 0 116032 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1028
timestamp 1669390400
transform 1 0 116480 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1031
timestamp 1669390400
transform 1 0 116816 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1095
timestamp 1669390400
transform 1 0 123984 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1099
timestamp 1669390400
transform 1 0 124432 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1102
timestamp 1669390400
transform 1 0 124768 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1166
timestamp 1669390400
transform 1 0 131936 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1170
timestamp 1669390400
transform 1 0 132384 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_1173
timestamp 1669390400
transform 1 0 132720 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_1237
timestamp 1669390400
transform 1 0 139888 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1241
timestamp 1669390400
transform 1 0 140336 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_1244
timestamp 1669390400
transform 1 0 140672 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_1276
timestamp 1669390400
transform 1 0 144256 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_1279
timestamp 1669390400
transform 1 0 144592 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_1295
timestamp 1669390400
transform 1 0 146384 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_1311
timestamp 1669390400
transform 1 0 148176 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1669390400
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1669390400
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_137
timestamp 1669390400
transform 1 0 16688 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_208
timestamp 1669390400
transform 1 0 24640 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_279
timestamp 1669390400
transform 1 0 32592 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1669390400
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1669390400
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_421
timestamp 1669390400
transform 1 0 48496 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1669390400
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_428
timestamp 1669390400
transform 1 0 49280 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_492
timestamp 1669390400
transform 1 0 56448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1669390400
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_499
timestamp 1669390400
transform 1 0 57232 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_563
timestamp 1669390400
transform 1 0 64400 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_567
timestamp 1669390400
transform 1 0 64848 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_570
timestamp 1669390400
transform 1 0 65184 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_634
timestamp 1669390400
transform 1 0 72352 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_638
timestamp 1669390400
transform 1 0 72800 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_641
timestamp 1669390400
transform 1 0 73136 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_705
timestamp 1669390400
transform 1 0 80304 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_709
timestamp 1669390400
transform 1 0 80752 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_712
timestamp 1669390400
transform 1 0 81088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_776
timestamp 1669390400
transform 1 0 88256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_780
timestamp 1669390400
transform 1 0 88704 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_783
timestamp 1669390400
transform 1 0 89040 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_847
timestamp 1669390400
transform 1 0 96208 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_851
timestamp 1669390400
transform 1 0 96656 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_854
timestamp 1669390400
transform 1 0 96992 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_918
timestamp 1669390400
transform 1 0 104160 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_922
timestamp 1669390400
transform 1 0 104608 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_925
timestamp 1669390400
transform 1 0 104944 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_989
timestamp 1669390400
transform 1 0 112112 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_993
timestamp 1669390400
transform 1 0 112560 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_996
timestamp 1669390400
transform 1 0 112896 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1060
timestamp 1669390400
transform 1 0 120064 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1064
timestamp 1669390400
transform 1 0 120512 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1067
timestamp 1669390400
transform 1 0 120848 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1131
timestamp 1669390400
transform 1 0 128016 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1135
timestamp 1669390400
transform 1 0 128464 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1138
timestamp 1669390400
transform 1 0 128800 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_1202
timestamp 1669390400
transform 1 0 135968 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1206
timestamp 1669390400
transform 1 0 136416 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_1209
timestamp 1669390400
transform 1 0 136752 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_1273
timestamp 1669390400
transform 1 0 143920 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1277
timestamp 1669390400
transform 1 0 144368 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_1280
timestamp 1669390400
transform 1 0 144704 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_1295
timestamp 1669390400
transform 1 0 146384 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_1311
timestamp 1669390400
transform 1 0 148176 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1669390400
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_172
timestamp 1669390400
transform 1 0 20608 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_243
timestamp 1669390400
transform 1 0 28560 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1669390400
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1669390400
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1669390400
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_456
timestamp 1669390400
transform 1 0 52416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1669390400
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_463
timestamp 1669390400
transform 1 0 53200 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_527
timestamp 1669390400
transform 1 0 60368 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_531
timestamp 1669390400
transform 1 0 60816 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_534
timestamp 1669390400
transform 1 0 61152 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_598
timestamp 1669390400
transform 1 0 68320 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_602
timestamp 1669390400
transform 1 0 68768 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_605
timestamp 1669390400
transform 1 0 69104 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_669
timestamp 1669390400
transform 1 0 76272 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_673
timestamp 1669390400
transform 1 0 76720 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_676
timestamp 1669390400
transform 1 0 77056 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_740
timestamp 1669390400
transform 1 0 84224 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_744
timestamp 1669390400
transform 1 0 84672 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_747
timestamp 1669390400
transform 1 0 85008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_811
timestamp 1669390400
transform 1 0 92176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_815
timestamp 1669390400
transform 1 0 92624 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_818
timestamp 1669390400
transform 1 0 92960 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_882
timestamp 1669390400
transform 1 0 100128 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_886
timestamp 1669390400
transform 1 0 100576 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_889
timestamp 1669390400
transform 1 0 100912 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_953
timestamp 1669390400
transform 1 0 108080 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_957
timestamp 1669390400
transform 1 0 108528 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_960
timestamp 1669390400
transform 1 0 108864 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1024
timestamp 1669390400
transform 1 0 116032 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1028
timestamp 1669390400
transform 1 0 116480 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1031
timestamp 1669390400
transform 1 0 116816 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1095
timestamp 1669390400
transform 1 0 123984 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1099
timestamp 1669390400
transform 1 0 124432 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1102
timestamp 1669390400
transform 1 0 124768 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1166
timestamp 1669390400
transform 1 0 131936 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1170
timestamp 1669390400
transform 1 0 132384 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_1173
timestamp 1669390400
transform 1 0 132720 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_1237
timestamp 1669390400
transform 1 0 139888 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1241
timestamp 1669390400
transform 1 0 140336 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_1244
timestamp 1669390400
transform 1 0 140672 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_1276
timestamp 1669390400
transform 1 0 144256 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_1279
timestamp 1669390400
transform 1 0 144592 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_1295
timestamp 1669390400
transform 1 0 146384 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_1311
timestamp 1669390400
transform 1 0 148176 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1669390400
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_137
timestamp 1669390400
transform 1 0 16688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1669390400
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_208
timestamp 1669390400
transform 1 0 24640 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1669390400
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_279
timestamp 1669390400
transform 1 0 32592 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1669390400
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1669390400
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_421
timestamp 1669390400
transform 1 0 48496 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_425
timestamp 1669390400
transform 1 0 48944 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_428
timestamp 1669390400
transform 1 0 49280 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_492
timestamp 1669390400
transform 1 0 56448 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_496
timestamp 1669390400
transform 1 0 56896 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_499
timestamp 1669390400
transform 1 0 57232 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_563
timestamp 1669390400
transform 1 0 64400 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_567
timestamp 1669390400
transform 1 0 64848 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_570
timestamp 1669390400
transform 1 0 65184 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_634
timestamp 1669390400
transform 1 0 72352 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_638
timestamp 1669390400
transform 1 0 72800 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_641
timestamp 1669390400
transform 1 0 73136 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_705
timestamp 1669390400
transform 1 0 80304 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_709
timestamp 1669390400
transform 1 0 80752 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_712
timestamp 1669390400
transform 1 0 81088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_776
timestamp 1669390400
transform 1 0 88256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_780
timestamp 1669390400
transform 1 0 88704 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_783
timestamp 1669390400
transform 1 0 89040 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_847
timestamp 1669390400
transform 1 0 96208 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_851
timestamp 1669390400
transform 1 0 96656 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_854
timestamp 1669390400
transform 1 0 96992 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_918
timestamp 1669390400
transform 1 0 104160 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_922
timestamp 1669390400
transform 1 0 104608 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_925
timestamp 1669390400
transform 1 0 104944 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_989
timestamp 1669390400
transform 1 0 112112 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_993
timestamp 1669390400
transform 1 0 112560 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_996
timestamp 1669390400
transform 1 0 112896 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1060
timestamp 1669390400
transform 1 0 120064 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1064
timestamp 1669390400
transform 1 0 120512 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1067
timestamp 1669390400
transform 1 0 120848 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1131
timestamp 1669390400
transform 1 0 128016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1135
timestamp 1669390400
transform 1 0 128464 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1138
timestamp 1669390400
transform 1 0 128800 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1202
timestamp 1669390400
transform 1 0 135968 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1206
timestamp 1669390400
transform 1 0 136416 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_1209
timestamp 1669390400
transform 1 0 136752 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_1273
timestamp 1669390400
transform 1 0 143920 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1277
timestamp 1669390400
transform 1 0 144368 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_1280
timestamp 1669390400
transform 1 0 144704 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_1312
timestamp 1669390400
transform 1 0 148288 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1669390400
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_101
timestamp 1669390400
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_172
timestamp 1669390400
transform 1 0 20608 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_243
timestamp 1669390400
transform 1 0 28560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_314
timestamp 1669390400
transform 1 0 36512 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1669390400
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1669390400
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_456
timestamp 1669390400
transform 1 0 52416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1669390400
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_463
timestamp 1669390400
transform 1 0 53200 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_527
timestamp 1669390400
transform 1 0 60368 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_531
timestamp 1669390400
transform 1 0 60816 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_534
timestamp 1669390400
transform 1 0 61152 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_598
timestamp 1669390400
transform 1 0 68320 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_602
timestamp 1669390400
transform 1 0 68768 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_605
timestamp 1669390400
transform 1 0 69104 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_669
timestamp 1669390400
transform 1 0 76272 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_673
timestamp 1669390400
transform 1 0 76720 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_676
timestamp 1669390400
transform 1 0 77056 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_740
timestamp 1669390400
transform 1 0 84224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_744
timestamp 1669390400
transform 1 0 84672 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_747
timestamp 1669390400
transform 1 0 85008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_811
timestamp 1669390400
transform 1 0 92176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_815
timestamp 1669390400
transform 1 0 92624 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_818
timestamp 1669390400
transform 1 0 92960 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_882
timestamp 1669390400
transform 1 0 100128 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_886
timestamp 1669390400
transform 1 0 100576 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_889
timestamp 1669390400
transform 1 0 100912 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_953
timestamp 1669390400
transform 1 0 108080 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_957
timestamp 1669390400
transform 1 0 108528 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_960
timestamp 1669390400
transform 1 0 108864 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1024
timestamp 1669390400
transform 1 0 116032 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1028
timestamp 1669390400
transform 1 0 116480 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1031
timestamp 1669390400
transform 1 0 116816 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1095
timestamp 1669390400
transform 1 0 123984 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1099
timestamp 1669390400
transform 1 0 124432 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1102
timestamp 1669390400
transform 1 0 124768 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1166
timestamp 1669390400
transform 1 0 131936 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1170
timestamp 1669390400
transform 1 0 132384 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_1173
timestamp 1669390400
transform 1 0 132720 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_1237
timestamp 1669390400
transform 1 0 139888 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1241
timestamp 1669390400
transform 1 0 140336 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_1244
timestamp 1669390400
transform 1 0 140672 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_1276
timestamp 1669390400
transform 1 0 144256 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1279
timestamp 1669390400
transform 1 0 144592 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_1295
timestamp 1669390400
transform 1 0 146384 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_1311
timestamp 1669390400
transform 1 0 148176 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1669390400
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1669390400
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_137
timestamp 1669390400
transform 1 0 16688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1669390400
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_208
timestamp 1669390400
transform 1 0 24640 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1669390400
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_279
timestamp 1669390400
transform 1 0 32592 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1669390400
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_421
timestamp 1669390400
transform 1 0 48496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1669390400
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_428
timestamp 1669390400
transform 1 0 49280 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_492
timestamp 1669390400
transform 1 0 56448 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1669390400
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_499
timestamp 1669390400
transform 1 0 57232 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_563
timestamp 1669390400
transform 1 0 64400 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_567
timestamp 1669390400
transform 1 0 64848 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_570
timestamp 1669390400
transform 1 0 65184 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_634
timestamp 1669390400
transform 1 0 72352 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_638
timestamp 1669390400
transform 1 0 72800 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_641
timestamp 1669390400
transform 1 0 73136 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_705
timestamp 1669390400
transform 1 0 80304 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_709
timestamp 1669390400
transform 1 0 80752 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_712
timestamp 1669390400
transform 1 0 81088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_776
timestamp 1669390400
transform 1 0 88256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_780
timestamp 1669390400
transform 1 0 88704 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_783
timestamp 1669390400
transform 1 0 89040 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_847
timestamp 1669390400
transform 1 0 96208 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_851
timestamp 1669390400
transform 1 0 96656 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_854
timestamp 1669390400
transform 1 0 96992 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_918
timestamp 1669390400
transform 1 0 104160 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_922
timestamp 1669390400
transform 1 0 104608 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_925
timestamp 1669390400
transform 1 0 104944 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_989
timestamp 1669390400
transform 1 0 112112 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_993
timestamp 1669390400
transform 1 0 112560 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_996
timestamp 1669390400
transform 1 0 112896 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1060
timestamp 1669390400
transform 1 0 120064 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1064
timestamp 1669390400
transform 1 0 120512 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_1067
timestamp 1669390400
transform 1 0 120848 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1131
timestamp 1669390400
transform 1 0 128016 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1135
timestamp 1669390400
transform 1 0 128464 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_1138
timestamp 1669390400
transform 1 0 128800 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_1202
timestamp 1669390400
transform 1 0 135968 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1206
timestamp 1669390400
transform 1 0 136416 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_1209
timestamp 1669390400
transform 1 0 136752 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1273
timestamp 1669390400
transform 1 0 143920 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1277
timestamp 1669390400
transform 1 0 144368 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_1280
timestamp 1669390400
transform 1 0 144704 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_1295
timestamp 1669390400
transform 1 0 146384 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_1311
timestamp 1669390400
transform 1 0 148176 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1669390400
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_101
timestamp 1669390400
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_172
timestamp 1669390400
transform 1 0 20608 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1669390400
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_314
timestamp 1669390400
transform 1 0 36512 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_318
timestamp 1669390400
transform 1 0 36960 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1669390400
transform 1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1669390400
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_456
timestamp 1669390400
transform 1 0 52416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1669390400
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_463
timestamp 1669390400
transform 1 0 53200 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_527
timestamp 1669390400
transform 1 0 60368 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_531
timestamp 1669390400
transform 1 0 60816 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_534
timestamp 1669390400
transform 1 0 61152 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_598
timestamp 1669390400
transform 1 0 68320 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_602
timestamp 1669390400
transform 1 0 68768 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_605
timestamp 1669390400
transform 1 0 69104 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_669
timestamp 1669390400
transform 1 0 76272 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_673
timestamp 1669390400
transform 1 0 76720 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_676
timestamp 1669390400
transform 1 0 77056 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_740
timestamp 1669390400
transform 1 0 84224 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_744
timestamp 1669390400
transform 1 0 84672 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_747
timestamp 1669390400
transform 1 0 85008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_811
timestamp 1669390400
transform 1 0 92176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_815
timestamp 1669390400
transform 1 0 92624 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_818
timestamp 1669390400
transform 1 0 92960 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_882
timestamp 1669390400
transform 1 0 100128 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_886
timestamp 1669390400
transform 1 0 100576 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_889
timestamp 1669390400
transform 1 0 100912 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_953
timestamp 1669390400
transform 1 0 108080 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_957
timestamp 1669390400
transform 1 0 108528 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_960
timestamp 1669390400
transform 1 0 108864 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1024
timestamp 1669390400
transform 1 0 116032 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1028
timestamp 1669390400
transform 1 0 116480 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_1031
timestamp 1669390400
transform 1 0 116816 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1095
timestamp 1669390400
transform 1 0 123984 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1099
timestamp 1669390400
transform 1 0 124432 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_1102
timestamp 1669390400
transform 1 0 124768 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1166
timestamp 1669390400
transform 1 0 131936 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1170
timestamp 1669390400
transform 1 0 132384 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_1173
timestamp 1669390400
transform 1 0 132720 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_1237
timestamp 1669390400
transform 1 0 139888 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1241
timestamp 1669390400
transform 1 0 140336 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_1244
timestamp 1669390400
transform 1 0 140672 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_1276
timestamp 1669390400
transform 1 0 144256 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1279
timestamp 1669390400
transform 1 0 144592 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1295
timestamp 1669390400
transform 1 0 146384 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1299
timestamp 1669390400
transform 1 0 146832 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_1303
timestamp 1669390400
transform 1 0 147280 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_1311
timestamp 1669390400
transform 1 0 148176 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_66
timestamp 1669390400
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1669390400
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_137
timestamp 1669390400
transform 1 0 16688 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_208
timestamp 1669390400
transform 1 0 24640 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_279
timestamp 1669390400
transform 1 0 32592 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1669390400
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_350
timestamp 1669390400
transform 1 0 40544 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_421
timestamp 1669390400
transform 1 0 48496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1669390400
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_428
timestamp 1669390400
transform 1 0 49280 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_492
timestamp 1669390400
transform 1 0 56448 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_496
timestamp 1669390400
transform 1 0 56896 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_499
timestamp 1669390400
transform 1 0 57232 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_563
timestamp 1669390400
transform 1 0 64400 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_567
timestamp 1669390400
transform 1 0 64848 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_570
timestamp 1669390400
transform 1 0 65184 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_634
timestamp 1669390400
transform 1 0 72352 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_638
timestamp 1669390400
transform 1 0 72800 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_641
timestamp 1669390400
transform 1 0 73136 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_705
timestamp 1669390400
transform 1 0 80304 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_709
timestamp 1669390400
transform 1 0 80752 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_712
timestamp 1669390400
transform 1 0 81088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_776
timestamp 1669390400
transform 1 0 88256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_780
timestamp 1669390400
transform 1 0 88704 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_783
timestamp 1669390400
transform 1 0 89040 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_847
timestamp 1669390400
transform 1 0 96208 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_851
timestamp 1669390400
transform 1 0 96656 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_854
timestamp 1669390400
transform 1 0 96992 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_918
timestamp 1669390400
transform 1 0 104160 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_922
timestamp 1669390400
transform 1 0 104608 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_925
timestamp 1669390400
transform 1 0 104944 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_989
timestamp 1669390400
transform 1 0 112112 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_993
timestamp 1669390400
transform 1 0 112560 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_996
timestamp 1669390400
transform 1 0 112896 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1060
timestamp 1669390400
transform 1 0 120064 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1064
timestamp 1669390400
transform 1 0 120512 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_1067
timestamp 1669390400
transform 1 0 120848 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1131
timestamp 1669390400
transform 1 0 128016 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1135
timestamp 1669390400
transform 1 0 128464 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_1138
timestamp 1669390400
transform 1 0 128800 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1202
timestamp 1669390400
transform 1 0 135968 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1206
timestamp 1669390400
transform 1 0 136416 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_1209
timestamp 1669390400
transform 1 0 136752 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_1241
timestamp 1669390400
transform 1 0 140336 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_1257
timestamp 1669390400
transform 1 0 142128 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_1265
timestamp 1669390400
transform 1 0 143024 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1269
timestamp 1669390400
transform 1 0 143472 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1273
timestamp 1669390400
transform 1 0 143920 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1277
timestamp 1669390400
transform 1 0 144368 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_1280
timestamp 1669390400
transform 1 0 144704 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1295
timestamp 1669390400
transform 1 0 146384 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_1311
timestamp 1669390400
transform 1 0 148176 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_69
timestamp 1669390400
transform 1 0 9072 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_72
timestamp 1669390400
transform 1 0 9408 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_104
timestamp 1669390400
transform 1 0 12992 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_107
timestamp 1669390400
transform 1 0 13328 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_139
timestamp 1669390400
transform 1 0 16912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_142
timestamp 1669390400
transform 1 0 17248 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_174
timestamp 1669390400
transform 1 0 20832 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_177
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_209
timestamp 1669390400
transform 1 0 24752 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_212
timestamp 1669390400
transform 1 0 25088 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_244
timestamp 1669390400
transform 1 0 28672 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_247
timestamp 1669390400
transform 1 0 29008 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_279
timestamp 1669390400
transform 1 0 32592 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_282
timestamp 1669390400
transform 1 0 32928 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_314
timestamp 1669390400
transform 1 0 36512 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_317
timestamp 1669390400
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_349
timestamp 1669390400
transform 1 0 40432 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_352
timestamp 1669390400
transform 1 0 40768 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_384
timestamp 1669390400
transform 1 0 44352 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_387
timestamp 1669390400
transform 1 0 44688 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_419
timestamp 1669390400
transform 1 0 48272 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_422
timestamp 1669390400
transform 1 0 48608 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_454
timestamp 1669390400
transform 1 0 52192 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_457
timestamp 1669390400
transform 1 0 52528 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_489
timestamp 1669390400
transform 1 0 56112 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_492
timestamp 1669390400
transform 1 0 56448 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_524
timestamp 1669390400
transform 1 0 60032 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_527
timestamp 1669390400
transform 1 0 60368 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_559
timestamp 1669390400
transform 1 0 63952 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_562
timestamp 1669390400
transform 1 0 64288 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_594
timestamp 1669390400
transform 1 0 67872 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_597
timestamp 1669390400
transform 1 0 68208 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_629
timestamp 1669390400
transform 1 0 71792 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_632
timestamp 1669390400
transform 1 0 72128 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_664
timestamp 1669390400
transform 1 0 75712 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_667
timestamp 1669390400
transform 1 0 76048 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_699
timestamp 1669390400
transform 1 0 79632 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_702
timestamp 1669390400
transform 1 0 79968 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_734
timestamp 1669390400
transform 1 0 83552 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_737
timestamp 1669390400
transform 1 0 83888 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_769
timestamp 1669390400
transform 1 0 87472 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_772
timestamp 1669390400
transform 1 0 87808 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_804
timestamp 1669390400
transform 1 0 91392 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_807
timestamp 1669390400
transform 1 0 91728 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_839
timestamp 1669390400
transform 1 0 95312 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_842
timestamp 1669390400
transform 1 0 95648 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_874
timestamp 1669390400
transform 1 0 99232 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_877
timestamp 1669390400
transform 1 0 99568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_909
timestamp 1669390400
transform 1 0 103152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_912
timestamp 1669390400
transform 1 0 103488 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_944
timestamp 1669390400
transform 1 0 107072 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_947
timestamp 1669390400
transform 1 0 107408 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_979
timestamp 1669390400
transform 1 0 110992 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_982
timestamp 1669390400
transform 1 0 111328 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1014
timestamp 1669390400
transform 1 0 114912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_1017
timestamp 1669390400
transform 1 0 115248 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1049
timestamp 1669390400
transform 1 0 118832 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_1052
timestamp 1669390400
transform 1 0 119168 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1084
timestamp 1669390400
transform 1 0 122752 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_1087
timestamp 1669390400
transform 1 0 123088 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1119
timestamp 1669390400
transform 1 0 126672 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_1122
timestamp 1669390400
transform 1 0 127008 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1154
timestamp 1669390400
transform 1 0 130592 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_1157
timestamp 1669390400
transform 1 0 130928 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1189
timestamp 1669390400
transform 1 0 134512 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_1192
timestamp 1669390400
transform 1 0 134848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1224
timestamp 1669390400
transform 1 0 138432 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_1227
timestamp 1669390400
transform 1 0 138768 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_1243
timestamp 1669390400
transform 1 0 140560 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_1251
timestamp 1669390400
transform 1 0 141456 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1255
timestamp 1669390400
transform 1 0 141904 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1259
timestamp 1669390400
transform 1 0 142352 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1262
timestamp 1669390400
transform 1 0 142688 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_1278
timestamp 1669390400
transform 1 0 144480 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1294
timestamp 1669390400
transform 1 0 146272 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1297
timestamp 1669390400
transform 1 0 146608 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_1312
timestamp 1669390400
transform 1 0 148288 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 148624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 148624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 148624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 148624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 148624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 148624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 148624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 148624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 148624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 148624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 148624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 148624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 148624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 148624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 148624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 148624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 148624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 148624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 148624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 148624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 148624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 148624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 148624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 148624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 148624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 148624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 148624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 148624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 148624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 148624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 148624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 148624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 148624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 148624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 148624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 148624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 148624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 148624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 148624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 148624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 148624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 148624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 148624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_86 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_87
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_88
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_89
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_90
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_91
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_92
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_93
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_94
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_95
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_96
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_97
timestamp 1669390400
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_98
timestamp 1669390400
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_99
timestamp 1669390400
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_100
timestamp 1669390400
transform 1 0 60144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_101
timestamp 1669390400
transform 1 0 64064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_102
timestamp 1669390400
transform 1 0 67984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_103
timestamp 1669390400
transform 1 0 71904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_104
timestamp 1669390400
transform 1 0 75824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_105
timestamp 1669390400
transform 1 0 79744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_106
timestamp 1669390400
transform 1 0 83664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_107
timestamp 1669390400
transform 1 0 87584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_108
timestamp 1669390400
transform 1 0 91504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_109
timestamp 1669390400
transform 1 0 95424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110
timestamp 1669390400
transform 1 0 99344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1669390400
transform 1 0 103264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1669390400
transform 1 0 107184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1669390400
transform 1 0 111104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1669390400
transform 1 0 115024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1669390400
transform 1 0 118944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1669390400
transform 1 0 122864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1669390400
transform 1 0 126784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1669390400
transform 1 0 130704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1669390400
transform 1 0 134624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1669390400
transform 1 0 138544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1669390400
transform 1 0 142464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1669390400
transform 1 0 146384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1669390400
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1669390400
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1669390400
transform 1 0 64960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1669390400
transform 1 0 72912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1669390400
transform 1 0 80864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1669390400
transform 1 0 88816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1669390400
transform 1 0 96768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1669390400
transform 1 0 104720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1669390400
transform 1 0 112672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1669390400
transform 1 0 120624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1669390400
transform 1 0 128576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1669390400
transform 1 0 136528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1669390400
transform 1 0 144480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1669390400
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1669390400
transform 1 0 60928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1669390400
transform 1 0 68880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1669390400
transform 1 0 76832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1669390400
transform 1 0 84784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1669390400
transform 1 0 92736 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1669390400
transform 1 0 100688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1669390400
transform 1 0 108640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1669390400
transform 1 0 116592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1669390400
transform 1 0 124544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1669390400
transform 1 0 132496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1669390400
transform 1 0 140448 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1669390400
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1669390400
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1669390400
transform 1 0 64960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1669390400
transform 1 0 72912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1669390400
transform 1 0 80864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1669390400
transform 1 0 88816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1669390400
transform 1 0 96768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1669390400
transform 1 0 104720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1669390400
transform 1 0 112672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1669390400
transform 1 0 120624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1669390400
transform 1 0 128576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1669390400
transform 1 0 136528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1669390400
transform 1 0 144480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1669390400
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1669390400
transform 1 0 60928 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1669390400
transform 1 0 68880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1669390400
transform 1 0 76832 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1669390400
transform 1 0 84784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1669390400
transform 1 0 92736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 100688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 108640 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 116592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 124544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 132496 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 140448 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 64960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 72912 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 80864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 88816 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 96768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 104720 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 112672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 120624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 128576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 136528 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 144480 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 60928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 68880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 76832 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 84784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 92736 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 100688 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 108640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 116592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 124544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 132496 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 140448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 64960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 72912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 80864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 88816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 96768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 104720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 112672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 120624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 128576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 136528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 144480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 60928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 68880 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 76832 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 84784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 92736 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 100688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 108640 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 116592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 124544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 132496 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 140448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 64960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 72912 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 80864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 88816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 96768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 104720 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 112672 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 120624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 128576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 136528 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 144480 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 60928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 68880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 76832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 84784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 92736 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 100688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 108640 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 116592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 124544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 132496 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 140448 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 64960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 72912 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 80864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 88816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 96768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 104720 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 112672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 120624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 128576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 136528 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 144480 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 60928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 68880 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 76832 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 84784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 92736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 100688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 108640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 116592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 124544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 132496 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 140448 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 64960 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 72912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 80864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 88816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 96768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 104720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 112672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 120624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 128576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 136528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 144480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 60928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 68880 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 76832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 84784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 92736 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 100688 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 108640 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 116592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 124544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 132496 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 140448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 64960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 72912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 80864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 88816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 96768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 104720 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 112672 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 120624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 128576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 136528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 144480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 60928 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 68880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 76832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 84784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 92736 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 100688 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 108640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 116592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 124544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 132496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 140448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 64960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 72912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 80864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 88816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 96768 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1669390400
transform 1 0 104720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1669390400
transform 1 0 112672 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1669390400
transform 1 0 120624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1669390400
transform 1 0 128576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1669390400
transform 1 0 136528 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1669390400
transform 1 0 144480 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1669390400
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1669390400
transform 1 0 60928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1669390400
transform 1 0 68880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1669390400
transform 1 0 76832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1669390400
transform 1 0 84784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1669390400
transform 1 0 92736 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1669390400
transform 1 0 100688 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1669390400
transform 1 0 108640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1669390400
transform 1 0 116592 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1669390400
transform 1 0 124544 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1669390400
transform 1 0 132496 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1669390400
transform 1 0 140448 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1669390400
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1669390400
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1669390400
transform 1 0 64960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1669390400
transform 1 0 72912 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1669390400
transform 1 0 80864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1669390400
transform 1 0 88816 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1669390400
transform 1 0 96768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1669390400
transform 1 0 104720 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1669390400
transform 1 0 112672 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1669390400
transform 1 0 120624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1669390400
transform 1 0 128576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1669390400
transform 1 0 136528 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1669390400
transform 1 0 144480 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1669390400
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1669390400
transform 1 0 60928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1669390400
transform 1 0 68880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1669390400
transform 1 0 76832 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1669390400
transform 1 0 84784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1669390400
transform 1 0 92736 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1669390400
transform 1 0 100688 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1669390400
transform 1 0 108640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1669390400
transform 1 0 116592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1669390400
transform 1 0 124544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1669390400
transform 1 0 132496 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1669390400
transform 1 0 140448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1669390400
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1669390400
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1669390400
transform 1 0 64960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1669390400
transform 1 0 72912 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1669390400
transform 1 0 80864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1669390400
transform 1 0 88816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1669390400
transform 1 0 96768 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1669390400
transform 1 0 104720 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1669390400
transform 1 0 112672 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1669390400
transform 1 0 120624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1669390400
transform 1 0 128576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1669390400
transform 1 0 136528 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1669390400
transform 1 0 144480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1669390400
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1669390400
transform 1 0 60928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1669390400
transform 1 0 68880 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1669390400
transform 1 0 76832 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1669390400
transform 1 0 84784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1669390400
transform 1 0 92736 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1669390400
transform 1 0 100688 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1669390400
transform 1 0 108640 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1669390400
transform 1 0 116592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1669390400
transform 1 0 124544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1669390400
transform 1 0 132496 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1669390400
transform 1 0 140448 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1669390400
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1669390400
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1669390400
transform 1 0 64960 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1669390400
transform 1 0 72912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1669390400
transform 1 0 80864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1669390400
transform 1 0 88816 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1669390400
transform 1 0 96768 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1669390400
transform 1 0 104720 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1669390400
transform 1 0 112672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1669390400
transform 1 0 120624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1669390400
transform 1 0 128576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1669390400
transform 1 0 136528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1669390400
transform 1 0 144480 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1669390400
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1669390400
transform 1 0 60928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1669390400
transform 1 0 68880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1669390400
transform 1 0 76832 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1669390400
transform 1 0 84784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1669390400
transform 1 0 92736 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1669390400
transform 1 0 100688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1669390400
transform 1 0 108640 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1669390400
transform 1 0 116592 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1669390400
transform 1 0 124544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1669390400
transform 1 0 132496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1669390400
transform 1 0 140448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1669390400
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1669390400
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1669390400
transform 1 0 64960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1669390400
transform 1 0 72912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1669390400
transform 1 0 80864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1669390400
transform 1 0 88816 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1669390400
transform 1 0 96768 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1669390400
transform 1 0 104720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1669390400
transform 1 0 112672 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1669390400
transform 1 0 120624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1669390400
transform 1 0 128576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1669390400
transform 1 0 136528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1669390400
transform 1 0 144480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1669390400
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1669390400
transform 1 0 60928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1669390400
transform 1 0 68880 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1669390400
transform 1 0 76832 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1669390400
transform 1 0 84784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1669390400
transform 1 0 92736 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1669390400
transform 1 0 100688 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1669390400
transform 1 0 108640 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1669390400
transform 1 0 116592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1669390400
transform 1 0 124544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1669390400
transform 1 0 132496 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1669390400
transform 1 0 140448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1669390400
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1669390400
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1669390400
transform 1 0 64960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1669390400
transform 1 0 72912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1669390400
transform 1 0 80864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1669390400
transform 1 0 88816 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1669390400
transform 1 0 96768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1669390400
transform 1 0 104720 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1669390400
transform 1 0 112672 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1669390400
transform 1 0 120624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1669390400
transform 1 0 128576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1669390400
transform 1 0 136528 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1669390400
transform 1 0 144480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1669390400
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1669390400
transform 1 0 60928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1669390400
transform 1 0 68880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1669390400
transform 1 0 76832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1669390400
transform 1 0 84784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1669390400
transform 1 0 92736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1669390400
transform 1 0 100688 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1669390400
transform 1 0 108640 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1669390400
transform 1 0 116592 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1669390400
transform 1 0 124544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1669390400
transform 1 0 132496 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_626
timestamp 1669390400
transform 1 0 140448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_627
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_628
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_629
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_630
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_631
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_632
timestamp 1669390400
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_633
timestamp 1669390400
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_634
timestamp 1669390400
transform 1 0 64960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_635
timestamp 1669390400
transform 1 0 72912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_636
timestamp 1669390400
transform 1 0 80864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_637
timestamp 1669390400
transform 1 0 88816 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_638
timestamp 1669390400
transform 1 0 96768 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_639
timestamp 1669390400
transform 1 0 104720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_640
timestamp 1669390400
transform 1 0 112672 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_641
timestamp 1669390400
transform 1 0 120624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_642
timestamp 1669390400
transform 1 0 128576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_643
timestamp 1669390400
transform 1 0 136528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_644
timestamp 1669390400
transform 1 0 144480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_645
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_646
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_647
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_648
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_649
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_650
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_651
timestamp 1669390400
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_652
timestamp 1669390400
transform 1 0 60928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_653
timestamp 1669390400
transform 1 0 68880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_654
timestamp 1669390400
transform 1 0 76832 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_655
timestamp 1669390400
transform 1 0 84784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_656
timestamp 1669390400
transform 1 0 92736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_657
timestamp 1669390400
transform 1 0 100688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_658
timestamp 1669390400
transform 1 0 108640 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_659
timestamp 1669390400
transform 1 0 116592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_660
timestamp 1669390400
transform 1 0 124544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_661
timestamp 1669390400
transform 1 0 132496 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_662
timestamp 1669390400
transform 1 0 140448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_663
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_664
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_665
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_666
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_667
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_668
timestamp 1669390400
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_669
timestamp 1669390400
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_670
timestamp 1669390400
transform 1 0 64960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_671
timestamp 1669390400
transform 1 0 72912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_672
timestamp 1669390400
transform 1 0 80864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_673
timestamp 1669390400
transform 1 0 88816 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_674
timestamp 1669390400
transform 1 0 96768 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_675
timestamp 1669390400
transform 1 0 104720 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_676
timestamp 1669390400
transform 1 0 112672 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_677
timestamp 1669390400
transform 1 0 120624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_678
timestamp 1669390400
transform 1 0 128576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_679
timestamp 1669390400
transform 1 0 136528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_680
timestamp 1669390400
transform 1 0 144480 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_681
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_682
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_683
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_684
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_685
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_686
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_687
timestamp 1669390400
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_688
timestamp 1669390400
transform 1 0 60928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_689
timestamp 1669390400
transform 1 0 68880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_690
timestamp 1669390400
transform 1 0 76832 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_691
timestamp 1669390400
transform 1 0 84784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_692
timestamp 1669390400
transform 1 0 92736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_693
timestamp 1669390400
transform 1 0 100688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_694
timestamp 1669390400
transform 1 0 108640 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_695
timestamp 1669390400
transform 1 0 116592 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_696
timestamp 1669390400
transform 1 0 124544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_697
timestamp 1669390400
transform 1 0 132496 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_698
timestamp 1669390400
transform 1 0 140448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_699
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_700
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_701
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_702
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_703
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_704
timestamp 1669390400
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_705
timestamp 1669390400
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_706
timestamp 1669390400
transform 1 0 64960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_707
timestamp 1669390400
transform 1 0 72912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_708
timestamp 1669390400
transform 1 0 80864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_709
timestamp 1669390400
transform 1 0 88816 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_710
timestamp 1669390400
transform 1 0 96768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_711
timestamp 1669390400
transform 1 0 104720 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_712
timestamp 1669390400
transform 1 0 112672 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_713
timestamp 1669390400
transform 1 0 120624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_714
timestamp 1669390400
transform 1 0 128576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_715
timestamp 1669390400
transform 1 0 136528 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_716
timestamp 1669390400
transform 1 0 144480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_717
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_718
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_719
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_720
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_721
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_722
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_723
timestamp 1669390400
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_724
timestamp 1669390400
transform 1 0 60928 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_725
timestamp 1669390400
transform 1 0 68880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_726
timestamp 1669390400
transform 1 0 76832 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_727
timestamp 1669390400
transform 1 0 84784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_728
timestamp 1669390400
transform 1 0 92736 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_729
timestamp 1669390400
transform 1 0 100688 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_730
timestamp 1669390400
transform 1 0 108640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_731
timestamp 1669390400
transform 1 0 116592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_732
timestamp 1669390400
transform 1 0 124544 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_733
timestamp 1669390400
transform 1 0 132496 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_734
timestamp 1669390400
transform 1 0 140448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_735
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_736
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_737
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_738
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_739
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_740
timestamp 1669390400
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_741
timestamp 1669390400
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_742
timestamp 1669390400
transform 1 0 64960 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_743
timestamp 1669390400
transform 1 0 72912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_744
timestamp 1669390400
transform 1 0 80864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_745
timestamp 1669390400
transform 1 0 88816 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_746
timestamp 1669390400
transform 1 0 96768 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_747
timestamp 1669390400
transform 1 0 104720 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_748
timestamp 1669390400
transform 1 0 112672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_749
timestamp 1669390400
transform 1 0 120624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_750
timestamp 1669390400
transform 1 0 128576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_751
timestamp 1669390400
transform 1 0 136528 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_752
timestamp 1669390400
transform 1 0 144480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_753
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_754
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_755
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_756
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_757
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_758
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_759
timestamp 1669390400
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_760
timestamp 1669390400
transform 1 0 60928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_761
timestamp 1669390400
transform 1 0 68880 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_762
timestamp 1669390400
transform 1 0 76832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_763
timestamp 1669390400
transform 1 0 84784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_764
timestamp 1669390400
transform 1 0 92736 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_765
timestamp 1669390400
transform 1 0 100688 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_766
timestamp 1669390400
transform 1 0 108640 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_767
timestamp 1669390400
transform 1 0 116592 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_768
timestamp 1669390400
transform 1 0 124544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_769
timestamp 1669390400
transform 1 0 132496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_770
timestamp 1669390400
transform 1 0 140448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_771
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_772
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_773
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_774
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_775
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_776
timestamp 1669390400
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_777
timestamp 1669390400
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_778
timestamp 1669390400
transform 1 0 64960 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_779
timestamp 1669390400
transform 1 0 72912 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_780
timestamp 1669390400
transform 1 0 80864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_781
timestamp 1669390400
transform 1 0 88816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_782
timestamp 1669390400
transform 1 0 96768 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_783
timestamp 1669390400
transform 1 0 104720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_784
timestamp 1669390400
transform 1 0 112672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_785
timestamp 1669390400
transform 1 0 120624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_786
timestamp 1669390400
transform 1 0 128576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_787
timestamp 1669390400
transform 1 0 136528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_788
timestamp 1669390400
transform 1 0 144480 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_789
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_790
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_791
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_792
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_793
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_794
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_795
timestamp 1669390400
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_796
timestamp 1669390400
transform 1 0 60928 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_797
timestamp 1669390400
transform 1 0 68880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_798
timestamp 1669390400
transform 1 0 76832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_799
timestamp 1669390400
transform 1 0 84784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_800
timestamp 1669390400
transform 1 0 92736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_801
timestamp 1669390400
transform 1 0 100688 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_802
timestamp 1669390400
transform 1 0 108640 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_803
timestamp 1669390400
transform 1 0 116592 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_804
timestamp 1669390400
transform 1 0 124544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_805
timestamp 1669390400
transform 1 0 132496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_806
timestamp 1669390400
transform 1 0 140448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_807
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_808
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_809
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_810
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_811
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_812
timestamp 1669390400
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_813
timestamp 1669390400
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_814
timestamp 1669390400
transform 1 0 64960 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_815
timestamp 1669390400
transform 1 0 72912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_816
timestamp 1669390400
transform 1 0 80864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_817
timestamp 1669390400
transform 1 0 88816 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_818
timestamp 1669390400
transform 1 0 96768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_819
timestamp 1669390400
transform 1 0 104720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_820
timestamp 1669390400
transform 1 0 112672 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_821
timestamp 1669390400
transform 1 0 120624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_822
timestamp 1669390400
transform 1 0 128576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_823
timestamp 1669390400
transform 1 0 136528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_824
timestamp 1669390400
transform 1 0 144480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_825
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_826
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_827
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_828
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_829
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_830
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_831
timestamp 1669390400
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_832
timestamp 1669390400
transform 1 0 60928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_833
timestamp 1669390400
transform 1 0 68880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_834
timestamp 1669390400
transform 1 0 76832 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_835
timestamp 1669390400
transform 1 0 84784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_836
timestamp 1669390400
transform 1 0 92736 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_837
timestamp 1669390400
transform 1 0 100688 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_838
timestamp 1669390400
transform 1 0 108640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_839
timestamp 1669390400
transform 1 0 116592 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_840
timestamp 1669390400
transform 1 0 124544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_841
timestamp 1669390400
transform 1 0 132496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_842
timestamp 1669390400
transform 1 0 140448 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_843
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_844
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_845
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_846
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_847
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_848
timestamp 1669390400
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_849
timestamp 1669390400
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_850
timestamp 1669390400
transform 1 0 64960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_851
timestamp 1669390400
transform 1 0 72912 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_852
timestamp 1669390400
transform 1 0 80864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_853
timestamp 1669390400
transform 1 0 88816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_854
timestamp 1669390400
transform 1 0 96768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_855
timestamp 1669390400
transform 1 0 104720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_856
timestamp 1669390400
transform 1 0 112672 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_857
timestamp 1669390400
transform 1 0 120624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_858
timestamp 1669390400
transform 1 0 128576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_859
timestamp 1669390400
transform 1 0 136528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_860
timestamp 1669390400
transform 1 0 144480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_861
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_862
timestamp 1669390400
transform 1 0 9184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_863
timestamp 1669390400
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_864
timestamp 1669390400
transform 1 0 17024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_865
timestamp 1669390400
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_866
timestamp 1669390400
transform 1 0 24864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_867
timestamp 1669390400
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_868
timestamp 1669390400
transform 1 0 32704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_869
timestamp 1669390400
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_870
timestamp 1669390400
transform 1 0 40544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_871
timestamp 1669390400
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_872
timestamp 1669390400
transform 1 0 48384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_873
timestamp 1669390400
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_874
timestamp 1669390400
transform 1 0 56224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_875
timestamp 1669390400
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_876
timestamp 1669390400
transform 1 0 64064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_877
timestamp 1669390400
transform 1 0 67984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_878
timestamp 1669390400
transform 1 0 71904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_879
timestamp 1669390400
transform 1 0 75824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_880
timestamp 1669390400
transform 1 0 79744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_881
timestamp 1669390400
transform 1 0 83664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_882
timestamp 1669390400
transform 1 0 87584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_883
timestamp 1669390400
transform 1 0 91504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_884
timestamp 1669390400
transform 1 0 95424 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_885
timestamp 1669390400
transform 1 0 99344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_886
timestamp 1669390400
transform 1 0 103264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_887
timestamp 1669390400
transform 1 0 107184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_888
timestamp 1669390400
transform 1 0 111104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_889
timestamp 1669390400
transform 1 0 115024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_890
timestamp 1669390400
transform 1 0 118944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_891
timestamp 1669390400
transform 1 0 122864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_892
timestamp 1669390400
transform 1 0 126784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_893
timestamp 1669390400
transform 1 0 130704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_894
timestamp 1669390400
transform 1 0 134624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_895
timestamp 1669390400
transform 1 0 138544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_896
timestamp 1669390400
transform 1 0 142464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_897
timestamp 1669390400
transform 1 0 146384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _042_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 131488 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _043_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 130592 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _044_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 123424 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _045_
timestamp 1669390400
transform 1 0 123648 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _046_
timestamp 1669390400
transform -1 0 124208 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _047_
timestamp 1669390400
transform 1 0 124432 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _048_
timestamp 1669390400
transform -1 0 126560 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _049_
timestamp 1669390400
transform 1 0 125552 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _050_
timestamp 1669390400
transform -1 0 128240 0 -1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _051_
timestamp 1669390400
transform 1 0 127456 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _052_
timestamp 1669390400
transform 1 0 133168 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _053_
timestamp 1669390400
transform -1 0 130032 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _054_
timestamp 1669390400
transform 1 0 130032 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _055_
timestamp 1669390400
transform -1 0 130816 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _056_
timestamp 1669390400
transform 1 0 130928 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _057_
timestamp 1669390400
transform -1 0 132048 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _058_
timestamp 1669390400
transform 1 0 132832 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _059_
timestamp 1669390400
transform -1 0 132944 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _060_
timestamp 1669390400
transform 1 0 134288 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _061_
timestamp 1669390400
transform 1 0 132832 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _062_
timestamp 1669390400
transform -1 0 135744 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _063_
timestamp 1669390400
transform 1 0 136864 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _064_
timestamp 1669390400
transform -1 0 137648 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _065_
timestamp 1669390400
transform 1 0 140784 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _066_
timestamp 1669390400
transform -1 0 139552 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _067_
timestamp 1669390400
transform 1 0 141680 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _068_
timestamp 1669390400
transform -1 0 142464 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _069_
timestamp 1669390400
transform 1 0 143696 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _070_
timestamp 1669390400
transform 1 0 133056 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _071_
timestamp 1669390400
transform -1 0 141456 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _072_
timestamp 1669390400
transform 1 0 139440 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _073_
timestamp 1669390400
transform -1 0 139552 0 1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _074_
timestamp 1669390400
transform 1 0 138544 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _075_
timestamp 1669390400
transform -1 0 139552 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _076_
timestamp 1669390400
transform 1 0 137760 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _077_
timestamp 1669390400
transform 1 0 105056 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _078_
timestamp 1669390400
transform 1 0 105056 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _079_
timestamp 1669390400
transform -1 0 129808 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _080_
timestamp 1669390400
transform -1 0 104496 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _081_
timestamp 1669390400
transform -1 0 96544 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _082_
timestamp 1669390400
transform 1 0 101024 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _083_
timestamp 1669390400
transform -1 0 98448 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _084_
timestamp 1669390400
transform 1 0 101024 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _085_
timestamp 1669390400
transform -1 0 98784 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _086_
timestamp 1669390400
transform 1 0 100016 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _087_
timestamp 1669390400
transform -1 0 100352 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _088_
timestamp 1669390400
transform 1 0 101024 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _089_
timestamp 1669390400
transform -1 0 106512 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _090_
timestamp 1669390400
transform -1 0 103264 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _091_
timestamp 1669390400
transform 1 0 103152 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _092_
timestamp 1669390400
transform -1 0 104048 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _093_
timestamp 1669390400
transform 1 0 104048 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _094_
timestamp 1669390400
transform -1 0 105168 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _095_
timestamp 1669390400
transform 1 0 105056 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _096_
timestamp 1669390400
transform -1 0 107072 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _097_
timestamp 1669390400
transform 1 0 107296 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _098_
timestamp 1669390400
transform -1 0 111216 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _099_
timestamp 1669390400
transform -1 0 110656 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _100_
timestamp 1669390400
transform 1 0 110208 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _101_
timestamp 1669390400
transform -1 0 111216 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _102_
timestamp 1669390400
transform 1 0 111104 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _103_
timestamp 1669390400
transform -1 0 112560 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _104_
timestamp 1669390400
transform 1 0 111552 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _105_
timestamp 1669390400
transform -1 0 114464 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _106_
timestamp 1669390400
transform 1 0 113008 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _107_
timestamp 1669390400
transform -1 0 118272 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _108_
timestamp 1669390400
transform -1 0 116480 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _109_
timestamp 1669390400
transform 1 0 116928 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _110_
timestamp 1669390400
transform -1 0 117376 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _111_
timestamp 1669390400
transform 1 0 118832 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _112_
timestamp 1669390400
transform -1 0 118608 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _113_
timestamp 1669390400
transform 1 0 119728 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _114_
timestamp 1669390400
transform -1 0 119392 0 -1 6272
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _115_
timestamp 1669390400
transform 1 0 119616 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _116_
timestamp 1669390400
transform -1 0 76160 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _117_
timestamp 1669390400
transform -1 0 78512 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _118_
timestamp 1669390400
transform -1 0 80304 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _119_
timestamp 1669390400
transform -1 0 81200 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _120_
timestamp 1669390400
transform -1 0 83552 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _121_
timestamp 1669390400
transform -1 0 86688 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _122_
timestamp 1669390400
transform -1 0 86912 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _123_
timestamp 1669390400
transform -1 0 87920 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _124_
timestamp 1669390400
transform -1 0 89600 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _125_
timestamp 1669390400
transform 1 0 76944 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _126_
timestamp 1669390400
transform 1 0 78736 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _127_
timestamp 1669390400
transform 1 0 81200 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _128_
timestamp 1669390400
transform 1 0 81984 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _129_
timestamp 1669390400
transform 1 0 84336 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _130_
timestamp 1669390400
transform 1 0 85344 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _131_
timestamp 1669390400
transform 1 0 87696 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _132_
timestamp 1669390400
transform 1 0 89152 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _133_
timestamp 1669390400
transform 1 0 90048 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _134_
timestamp 1669390400
transform -1 0 73696 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _135_
timestamp 1669390400
transform 1 0 75264 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 146608 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input2
timestamp 1669390400
transform -1 0 144592 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform -1 0 146608 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input4
timestamp 1669390400
transform -1 0 146608 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input5
timestamp 1669390400
transform -1 0 146608 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input6
timestamp 1669390400
transform -1 0 146608 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input7
timestamp 1669390400
transform -1 0 146608 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input8
timestamp 1669390400
transform -1 0 146608 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input9
timestamp 1669390400
transform -1 0 146608 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input10
timestamp 1669390400
transform -1 0 146608 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input11
timestamp 1669390400
transform -1 0 144368 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input12
timestamp 1669390400
transform 1 0 22064 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input13
timestamp 1669390400
transform 1 0 38640 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input14
timestamp 1669390400
transform 1 0 41440 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input15
timestamp 1669390400
transform 1 0 42224 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input16
timestamp 1669390400
transform 1 0 43568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input17
timestamp 1669390400
transform 1 0 45584 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input18
timestamp 1669390400
transform 1 0 46480 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input19
timestamp 1669390400
transform 1 0 49392 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input20
timestamp 1669390400
transform 1 0 50400 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input21
timestamp 1669390400
transform 1 0 52304 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input22
timestamp 1669390400
transform 1 0 53984 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input23
timestamp 1669390400
transform 1 0 22960 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input24
timestamp 1669390400
transform 1 0 55104 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input25
timestamp 1669390400
transform 1 0 57344 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input26
timestamp 1669390400
transform 1 0 58240 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input27
timestamp 1669390400
transform 1 0 60704 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input28
timestamp 1669390400
transform 1 0 62160 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input29
timestamp 1669390400
transform 1 0 64064 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input30
timestamp 1669390400
transform 1 0 65744 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input31
timestamp 1669390400
transform 1 0 67088 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input32
timestamp 1669390400
transform 1 0 69104 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input33
timestamp 1669390400
transform 1 0 70000 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input34
timestamp 1669390400
transform 1 0 25536 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input35
timestamp 1669390400
transform 1 0 73248 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input36
timestamp 1669390400
transform 1 0 73920 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input37
timestamp 1669390400
transform 1 0 26880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input38
timestamp 1669390400
transform 1 0 28448 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input39
timestamp 1669390400
transform 1 0 30464 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input40
timestamp 1669390400
transform 1 0 30800 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input41
timestamp 1669390400
transform 1 0 33824 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input42
timestamp 1669390400
transform 1 0 34720 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input43
timestamp 1669390400
transform 1 0 37184 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input44
timestamp 1669390400
transform 1 0 92624 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input45
timestamp 1669390400
transform -1 0 111552 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input46
timestamp 1669390400
transform -1 0 113232 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input47
timestamp 1669390400
transform 1 0 113008 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input48
timestamp 1669390400
transform 1 0 115360 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input49
timestamp 1669390400
transform 1 0 116144 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input50
timestamp 1669390400
transform -1 0 119952 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input51
timestamp 1669390400
transform -1 0 121296 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input52
timestamp 1669390400
transform 1 0 121184 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input53
timestamp 1669390400
transform -1 0 124992 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input54
timestamp 1669390400
transform 1 0 124544 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input55
timestamp 1669390400
transform 1 0 94304 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input56
timestamp 1669390400
transform 1 0 127120 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input57
timestamp 1669390400
transform 1 0 128912 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input58
timestamp 1669390400
transform -1 0 132832 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input59
timestamp 1669390400
transform -1 0 133056 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input60
timestamp 1669390400
transform -1 0 135072 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input61
timestamp 1669390400
transform -1 0 136752 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input62
timestamp 1669390400
transform -1 0 138656 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input63
timestamp 1669390400
transform -1 0 140672 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input64
timestamp 1669390400
transform 1 0 139664 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input65
timestamp 1669390400
transform -1 0 143472 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input66
timestamp 1669390400
transform 1 0 95984 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input67
timestamp 1669390400
transform -1 0 144816 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input68
timestamp 1669390400
transform -1 0 144592 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input69
timestamp 1669390400
transform 1 0 97664 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input70
timestamp 1669390400
transform -1 0 101472 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input71
timestamp 1669390400
transform 1 0 101024 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input72
timestamp 1669390400
transform -1 0 105392 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input73
timestamp 1669390400
transform -1 0 106848 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input74
timestamp 1669390400
transform -1 0 109312 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input75
timestamp 1669390400
transform 1 0 107744 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output76 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 8512 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output77
timestamp 1669390400
transform -1 0 9072 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output78
timestamp 1669390400
transform -1 0 11200 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output79
timestamp 1669390400
transform -1 0 12992 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output80
timestamp 1669390400
transform -1 0 15120 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output81
timestamp 1669390400
transform -1 0 16912 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output82
timestamp 1669390400
transform -1 0 18928 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output83
timestamp 1669390400
transform -1 0 20272 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output84
timestamp 1669390400
transform -1 0 20832 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output85
timestamp 1669390400
transform 1 0 77952 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output86
timestamp 1669390400
transform 1 0 80080 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output87
timestamp 1669390400
transform 1 0 81872 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output88
timestamp 1669390400
transform 1 0 82544 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output89
timestamp 1669390400
transform -1 0 85792 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output90
timestamp 1669390400
transform 1 0 85904 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output91
timestamp 1669390400
transform 1 0 87920 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output92
timestamp 1669390400
transform 1 0 89712 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output93
timestamp 1669390400
transform 1 0 90944 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output94
timestamp 1669390400
transform -1 0 7168 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output95
timestamp 1669390400
transform 1 0 76160 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output96
timestamp 1669390400
transform 1 0 144816 0 1 10976
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output97
timestamp 1669390400
transform 1 0 144816 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output98
timestamp 1669390400
transform 1 0 144816 0 -1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output99
timestamp 1669390400
transform 1 0 144816 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output100
timestamp 1669390400
transform 1 0 144816 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output101
timestamp 1669390400
transform 1 0 144816 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output102
timestamp 1669390400
transform 1 0 144816 0 -1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output103
timestamp 1669390400
transform 1 0 144816 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output104
timestamp 1669390400
transform 1 0 144816 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output105
timestamp 1669390400
transform 1 0 144816 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output106
timestamp 1669390400
transform 1 0 144816 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output107
timestamp 1669390400
transform 1 0 144816 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output108
timestamp 1669390400
transform 1 0 144816 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output109
timestamp 1669390400
transform 1 0 144816 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output110
timestamp 1669390400
transform 1 0 144816 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output111
timestamp 1669390400
transform 1 0 144816 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output112
timestamp 1669390400
transform 1 0 144816 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output113
timestamp 1669390400
transform 1 0 144816 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output114
timestamp 1669390400
transform 1 0 144816 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output115
timestamp 1669390400
transform 1 0 144816 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output116
timestamp 1669390400
transform 1 0 144704 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output117
timestamp 1669390400
transform 1 0 146720 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output118
timestamp 1669390400
transform 1 0 144816 0 1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output119
timestamp 1669390400
transform 1 0 142912 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output120
timestamp 1669390400
transform 1 0 146608 0 -1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output121
timestamp 1669390400
transform 1 0 144816 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output122
timestamp 1669390400
transform 1 0 144816 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output123
timestamp 1669390400
transform 1 0 144816 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output124
timestamp 1669390400
transform 1 0 144816 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output125
timestamp 1669390400
transform 1 0 144816 0 1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output126
timestamp 1669390400
transform 1 0 144816 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output127
timestamp 1669390400
transform 1 0 144816 0 1 18816
box -86 -86 1654 870
<< labels >>
flabel metal3 s 149200 2016 150000 2128 0 FreeSans 448 0 0 0 addr[0]
port 0 nsew signal input
flabel metal3 s 149200 2912 150000 3024 0 FreeSans 448 0 0 0 addr[1]
port 1 nsew signal input
flabel metal3 s 149200 3808 150000 3920 0 FreeSans 448 0 0 0 addr[2]
port 2 nsew signal input
flabel metal3 s 149200 4704 150000 4816 0 FreeSans 448 0 0 0 addr[3]
port 3 nsew signal input
flabel metal3 s 149200 5600 150000 5712 0 FreeSans 448 0 0 0 addr[4]
port 4 nsew signal input
flabel metal3 s 149200 6496 150000 6608 0 FreeSans 448 0 0 0 addr[5]
port 5 nsew signal input
flabel metal3 s 149200 7392 150000 7504 0 FreeSans 448 0 0 0 addr[6]
port 6 nsew signal input
flabel metal3 s 149200 8288 150000 8400 0 FreeSans 448 0 0 0 addr[7]
port 7 nsew signal input
flabel metal3 s 149200 9184 150000 9296 0 FreeSans 448 0 0 0 addr[8]
port 8 nsew signal input
flabel metal3 s 149200 10080 150000 10192 0 FreeSans 448 0 0 0 addr[9]
port 9 nsew signal input
flabel metal2 s 6832 0 6944 800 0 FreeSans 448 90 0 0 addr_mem0[0]
port 10 nsew signal tristate
flabel metal2 s 8512 0 8624 800 0 FreeSans 448 90 0 0 addr_mem0[1]
port 11 nsew signal tristate
flabel metal2 s 10192 0 10304 800 0 FreeSans 448 90 0 0 addr_mem0[2]
port 12 nsew signal tristate
flabel metal2 s 11872 0 11984 800 0 FreeSans 448 90 0 0 addr_mem0[3]
port 13 nsew signal tristate
flabel metal2 s 13552 0 13664 800 0 FreeSans 448 90 0 0 addr_mem0[4]
port 14 nsew signal tristate
flabel metal2 s 15232 0 15344 800 0 FreeSans 448 90 0 0 addr_mem0[5]
port 15 nsew signal tristate
flabel metal2 s 16912 0 17024 800 0 FreeSans 448 90 0 0 addr_mem0[6]
port 16 nsew signal tristate
flabel metal2 s 18592 0 18704 800 0 FreeSans 448 90 0 0 addr_mem0[7]
port 17 nsew signal tristate
flabel metal2 s 20272 0 20384 800 0 FreeSans 448 90 0 0 addr_mem0[8]
port 18 nsew signal tristate
flabel metal2 s 77392 0 77504 800 0 FreeSans 448 90 0 0 addr_mem1[0]
port 19 nsew signal tristate
flabel metal2 s 79072 0 79184 800 0 FreeSans 448 90 0 0 addr_mem1[1]
port 20 nsew signal tristate
flabel metal2 s 80752 0 80864 800 0 FreeSans 448 90 0 0 addr_mem1[2]
port 21 nsew signal tristate
flabel metal2 s 82432 0 82544 800 0 FreeSans 448 90 0 0 addr_mem1[3]
port 22 nsew signal tristate
flabel metal2 s 84112 0 84224 800 0 FreeSans 448 90 0 0 addr_mem1[4]
port 23 nsew signal tristate
flabel metal2 s 85792 0 85904 800 0 FreeSans 448 90 0 0 addr_mem1[5]
port 24 nsew signal tristate
flabel metal2 s 87472 0 87584 800 0 FreeSans 448 90 0 0 addr_mem1[6]
port 25 nsew signal tristate
flabel metal2 s 89152 0 89264 800 0 FreeSans 448 90 0 0 addr_mem1[7]
port 26 nsew signal tristate
flabel metal2 s 90832 0 90944 800 0 FreeSans 448 90 0 0 addr_mem1[8]
port 27 nsew signal tristate
flabel metal3 s 149200 1120 150000 1232 0 FreeSans 448 0 0 0 csb
port 28 nsew signal input
flabel metal2 s 5152 0 5264 800 0 FreeSans 448 90 0 0 csb_mem0
port 29 nsew signal tristate
flabel metal2 s 75712 0 75824 800 0 FreeSans 448 90 0 0 csb_mem1
port 30 nsew signal tristate
flabel metal3 s 149200 10976 150000 11088 0 FreeSans 448 0 0 0 dout[0]
port 31 nsew signal tristate
flabel metal3 s 149200 19936 150000 20048 0 FreeSans 448 0 0 0 dout[10]
port 32 nsew signal tristate
flabel metal3 s 149200 20832 150000 20944 0 FreeSans 448 0 0 0 dout[11]
port 33 nsew signal tristate
flabel metal3 s 149200 21728 150000 21840 0 FreeSans 448 0 0 0 dout[12]
port 34 nsew signal tristate
flabel metal3 s 149200 22624 150000 22736 0 FreeSans 448 0 0 0 dout[13]
port 35 nsew signal tristate
flabel metal3 s 149200 23520 150000 23632 0 FreeSans 448 0 0 0 dout[14]
port 36 nsew signal tristate
flabel metal3 s 149200 24416 150000 24528 0 FreeSans 448 0 0 0 dout[15]
port 37 nsew signal tristate
flabel metal3 s 149200 25312 150000 25424 0 FreeSans 448 0 0 0 dout[16]
port 38 nsew signal tristate
flabel metal3 s 149200 26208 150000 26320 0 FreeSans 448 0 0 0 dout[17]
port 39 nsew signal tristate
flabel metal3 s 149200 27104 150000 27216 0 FreeSans 448 0 0 0 dout[18]
port 40 nsew signal tristate
flabel metal3 s 149200 28000 150000 28112 0 FreeSans 448 0 0 0 dout[19]
port 41 nsew signal tristate
flabel metal3 s 149200 11872 150000 11984 0 FreeSans 448 0 0 0 dout[1]
port 42 nsew signal tristate
flabel metal3 s 149200 28896 150000 29008 0 FreeSans 448 0 0 0 dout[20]
port 43 nsew signal tristate
flabel metal3 s 149200 29792 150000 29904 0 FreeSans 448 0 0 0 dout[21]
port 44 nsew signal tristate
flabel metal3 s 149200 30688 150000 30800 0 FreeSans 448 0 0 0 dout[22]
port 45 nsew signal tristate
flabel metal3 s 149200 31584 150000 31696 0 FreeSans 448 0 0 0 dout[23]
port 46 nsew signal tristate
flabel metal3 s 149200 32480 150000 32592 0 FreeSans 448 0 0 0 dout[24]
port 47 nsew signal tristate
flabel metal3 s 149200 33376 150000 33488 0 FreeSans 448 0 0 0 dout[25]
port 48 nsew signal tristate
flabel metal3 s 149200 34272 150000 34384 0 FreeSans 448 0 0 0 dout[26]
port 49 nsew signal tristate
flabel metal3 s 149200 35168 150000 35280 0 FreeSans 448 0 0 0 dout[27]
port 50 nsew signal tristate
flabel metal3 s 149200 36064 150000 36176 0 FreeSans 448 0 0 0 dout[28]
port 51 nsew signal tristate
flabel metal3 s 149200 36960 150000 37072 0 FreeSans 448 0 0 0 dout[29]
port 52 nsew signal tristate
flabel metal3 s 149200 12768 150000 12880 0 FreeSans 448 0 0 0 dout[2]
port 53 nsew signal tristate
flabel metal3 s 149200 37856 150000 37968 0 FreeSans 448 0 0 0 dout[30]
port 54 nsew signal tristate
flabel metal3 s 149200 38752 150000 38864 0 FreeSans 448 0 0 0 dout[31]
port 55 nsew signal tristate
flabel metal3 s 149200 13664 150000 13776 0 FreeSans 448 0 0 0 dout[3]
port 56 nsew signal tristate
flabel metal3 s 149200 14560 150000 14672 0 FreeSans 448 0 0 0 dout[4]
port 57 nsew signal tristate
flabel metal3 s 149200 15456 150000 15568 0 FreeSans 448 0 0 0 dout[5]
port 58 nsew signal tristate
flabel metal3 s 149200 16352 150000 16464 0 FreeSans 448 0 0 0 dout[6]
port 59 nsew signal tristate
flabel metal3 s 149200 17248 150000 17360 0 FreeSans 448 0 0 0 dout[7]
port 60 nsew signal tristate
flabel metal3 s 149200 18144 150000 18256 0 FreeSans 448 0 0 0 dout[8]
port 61 nsew signal tristate
flabel metal3 s 149200 19040 150000 19152 0 FreeSans 448 0 0 0 dout[9]
port 62 nsew signal tristate
flabel metal2 s 21952 0 22064 800 0 FreeSans 448 90 0 0 dout_mem0[0]
port 63 nsew signal input
flabel metal2 s 38752 0 38864 800 0 FreeSans 448 90 0 0 dout_mem0[10]
port 64 nsew signal input
flabel metal2 s 40432 0 40544 800 0 FreeSans 448 90 0 0 dout_mem0[11]
port 65 nsew signal input
flabel metal2 s 42112 0 42224 800 0 FreeSans 448 90 0 0 dout_mem0[12]
port 66 nsew signal input
flabel metal2 s 43792 0 43904 800 0 FreeSans 448 90 0 0 dout_mem0[13]
port 67 nsew signal input
flabel metal2 s 45472 0 45584 800 0 FreeSans 448 90 0 0 dout_mem0[14]
port 68 nsew signal input
flabel metal2 s 47152 0 47264 800 0 FreeSans 448 90 0 0 dout_mem0[15]
port 69 nsew signal input
flabel metal2 s 48832 0 48944 800 0 FreeSans 448 90 0 0 dout_mem0[16]
port 70 nsew signal input
flabel metal2 s 50512 0 50624 800 0 FreeSans 448 90 0 0 dout_mem0[17]
port 71 nsew signal input
flabel metal2 s 52192 0 52304 800 0 FreeSans 448 90 0 0 dout_mem0[18]
port 72 nsew signal input
flabel metal2 s 53872 0 53984 800 0 FreeSans 448 90 0 0 dout_mem0[19]
port 73 nsew signal input
flabel metal2 s 23632 0 23744 800 0 FreeSans 448 90 0 0 dout_mem0[1]
port 74 nsew signal input
flabel metal2 s 55552 0 55664 800 0 FreeSans 448 90 0 0 dout_mem0[20]
port 75 nsew signal input
flabel metal2 s 57232 0 57344 800 0 FreeSans 448 90 0 0 dout_mem0[21]
port 76 nsew signal input
flabel metal2 s 58912 0 59024 800 0 FreeSans 448 90 0 0 dout_mem0[22]
port 77 nsew signal input
flabel metal2 s 60592 0 60704 800 0 FreeSans 448 90 0 0 dout_mem0[23]
port 78 nsew signal input
flabel metal2 s 62272 0 62384 800 0 FreeSans 448 90 0 0 dout_mem0[24]
port 79 nsew signal input
flabel metal2 s 63952 0 64064 800 0 FreeSans 448 90 0 0 dout_mem0[25]
port 80 nsew signal input
flabel metal2 s 65632 0 65744 800 0 FreeSans 448 90 0 0 dout_mem0[26]
port 81 nsew signal input
flabel metal2 s 67312 0 67424 800 0 FreeSans 448 90 0 0 dout_mem0[27]
port 82 nsew signal input
flabel metal2 s 68992 0 69104 800 0 FreeSans 448 90 0 0 dout_mem0[28]
port 83 nsew signal input
flabel metal2 s 70672 0 70784 800 0 FreeSans 448 90 0 0 dout_mem0[29]
port 84 nsew signal input
flabel metal2 s 25312 0 25424 800 0 FreeSans 448 90 0 0 dout_mem0[2]
port 85 nsew signal input
flabel metal2 s 72352 0 72464 800 0 FreeSans 448 90 0 0 dout_mem0[30]
port 86 nsew signal input
flabel metal2 s 74032 0 74144 800 0 FreeSans 448 90 0 0 dout_mem0[31]
port 87 nsew signal input
flabel metal2 s 26992 0 27104 800 0 FreeSans 448 90 0 0 dout_mem0[3]
port 88 nsew signal input
flabel metal2 s 28672 0 28784 800 0 FreeSans 448 90 0 0 dout_mem0[4]
port 89 nsew signal input
flabel metal2 s 30352 0 30464 800 0 FreeSans 448 90 0 0 dout_mem0[5]
port 90 nsew signal input
flabel metal2 s 32032 0 32144 800 0 FreeSans 448 90 0 0 dout_mem0[6]
port 91 nsew signal input
flabel metal2 s 33712 0 33824 800 0 FreeSans 448 90 0 0 dout_mem0[7]
port 92 nsew signal input
flabel metal2 s 35392 0 35504 800 0 FreeSans 448 90 0 0 dout_mem0[8]
port 93 nsew signal input
flabel metal2 s 37072 0 37184 800 0 FreeSans 448 90 0 0 dout_mem0[9]
port 94 nsew signal input
flabel metal2 s 92512 0 92624 800 0 FreeSans 448 90 0 0 dout_mem1[0]
port 95 nsew signal input
flabel metal2 s 109312 0 109424 800 0 FreeSans 448 90 0 0 dout_mem1[10]
port 96 nsew signal input
flabel metal2 s 110992 0 111104 800 0 FreeSans 448 90 0 0 dout_mem1[11]
port 97 nsew signal input
flabel metal2 s 112672 0 112784 800 0 FreeSans 448 90 0 0 dout_mem1[12]
port 98 nsew signal input
flabel metal2 s 114352 0 114464 800 0 FreeSans 448 90 0 0 dout_mem1[13]
port 99 nsew signal input
flabel metal2 s 116032 0 116144 800 0 FreeSans 448 90 0 0 dout_mem1[14]
port 100 nsew signal input
flabel metal2 s 117712 0 117824 800 0 FreeSans 448 90 0 0 dout_mem1[15]
port 101 nsew signal input
flabel metal2 s 119392 0 119504 800 0 FreeSans 448 90 0 0 dout_mem1[16]
port 102 nsew signal input
flabel metal2 s 121072 0 121184 800 0 FreeSans 448 90 0 0 dout_mem1[17]
port 103 nsew signal input
flabel metal2 s 122752 0 122864 800 0 FreeSans 448 90 0 0 dout_mem1[18]
port 104 nsew signal input
flabel metal2 s 124432 0 124544 800 0 FreeSans 448 90 0 0 dout_mem1[19]
port 105 nsew signal input
flabel metal2 s 94192 0 94304 800 0 FreeSans 448 90 0 0 dout_mem1[1]
port 106 nsew signal input
flabel metal2 s 126112 0 126224 800 0 FreeSans 448 90 0 0 dout_mem1[20]
port 107 nsew signal input
flabel metal2 s 127792 0 127904 800 0 FreeSans 448 90 0 0 dout_mem1[21]
port 108 nsew signal input
flabel metal2 s 129472 0 129584 800 0 FreeSans 448 90 0 0 dout_mem1[22]
port 109 nsew signal input
flabel metal2 s 131152 0 131264 800 0 FreeSans 448 90 0 0 dout_mem1[23]
port 110 nsew signal input
flabel metal2 s 132832 0 132944 800 0 FreeSans 448 90 0 0 dout_mem1[24]
port 111 nsew signal input
flabel metal2 s 134512 0 134624 800 0 FreeSans 448 90 0 0 dout_mem1[25]
port 112 nsew signal input
flabel metal2 s 136192 0 136304 800 0 FreeSans 448 90 0 0 dout_mem1[26]
port 113 nsew signal input
flabel metal2 s 137872 0 137984 800 0 FreeSans 448 90 0 0 dout_mem1[27]
port 114 nsew signal input
flabel metal2 s 139552 0 139664 800 0 FreeSans 448 90 0 0 dout_mem1[28]
port 115 nsew signal input
flabel metal2 s 141232 0 141344 800 0 FreeSans 448 90 0 0 dout_mem1[29]
port 116 nsew signal input
flabel metal2 s 95872 0 95984 800 0 FreeSans 448 90 0 0 dout_mem1[2]
port 117 nsew signal input
flabel metal2 s 142912 0 143024 800 0 FreeSans 448 90 0 0 dout_mem1[30]
port 118 nsew signal input
flabel metal2 s 144592 0 144704 800 0 FreeSans 448 90 0 0 dout_mem1[31]
port 119 nsew signal input
flabel metal2 s 97552 0 97664 800 0 FreeSans 448 90 0 0 dout_mem1[3]
port 120 nsew signal input
flabel metal2 s 99232 0 99344 800 0 FreeSans 448 90 0 0 dout_mem1[4]
port 121 nsew signal input
flabel metal2 s 100912 0 101024 800 0 FreeSans 448 90 0 0 dout_mem1[5]
port 122 nsew signal input
flabel metal2 s 102592 0 102704 800 0 FreeSans 448 90 0 0 dout_mem1[6]
port 123 nsew signal input
flabel metal2 s 104272 0 104384 800 0 FreeSans 448 90 0 0 dout_mem1[7]
port 124 nsew signal input
flabel metal2 s 105952 0 106064 800 0 FreeSans 448 90 0 0 dout_mem1[8]
port 125 nsew signal input
flabel metal2 s 107632 0 107744 800 0 FreeSans 448 90 0 0 dout_mem1[9]
port 126 nsew signal input
flabel metal4 s 19594 3076 19914 36908 0 FreeSans 1280 90 0 0 vdd
port 127 nsew power bidirectional
flabel metal4 s 56414 3076 56734 36908 0 FreeSans 1280 90 0 0 vdd
port 127 nsew power bidirectional
flabel metal4 s 93234 3076 93554 36908 0 FreeSans 1280 90 0 0 vdd
port 127 nsew power bidirectional
flabel metal4 s 130054 3076 130374 36908 0 FreeSans 1280 90 0 0 vdd
port 127 nsew power bidirectional
flabel metal4 s 38004 3076 38324 36908 0 FreeSans 1280 90 0 0 vss
port 128 nsew ground bidirectional
flabel metal4 s 74824 3076 75144 36908 0 FreeSans 1280 90 0 0 vss
port 128 nsew ground bidirectional
flabel metal4 s 111644 3076 111964 36908 0 FreeSans 1280 90 0 0 vss
port 128 nsew ground bidirectional
flabel metal4 s 148464 3076 148784 36908 0 FreeSans 1280 90 0 0 vss
port 128 nsew ground bidirectional
rlabel metal1 74984 36848 74984 36848 0 vdd
rlabel via1 75064 36064 75064 36064 0 vss
rlabel metal3 123480 4984 123480 4984 0 _000_
rlabel metal3 124264 5880 124264 5880 0 _001_
rlabel metal2 126280 5600 126280 5600 0 _002_
rlabel metal2 127960 4592 127960 4592 0 _003_
rlabel metal2 132104 5880 132104 5880 0 _004_
rlabel metal2 129752 5936 129752 5936 0 _005_
rlabel metal3 130816 6104 130816 6104 0 _006_
rlabel metal3 132384 5320 132384 5320 0 _007_
rlabel metal3 133560 5880 133560 5880 0 _008_
rlabel metal3 139832 5096 139832 5096 0 _009_
rlabel metal3 136248 5320 136248 5320 0 _010_
rlabel metal2 140952 5992 140952 5992 0 _011_
rlabel metal3 140560 5320 140560 5320 0 _012_
rlabel metal3 143024 4424 143024 4424 0 _013_
rlabel metal2 140392 6608 140392 6608 0 _014_
rlabel metal3 140448 6104 140448 6104 0 _015_
rlabel metal2 139272 7168 139272 7168 0 _016_
rlabel metal2 137928 4424 137928 4424 0 _017_
rlabel metal2 105336 6776 105336 6776 0 _018_
rlabel metal2 118104 3696 118104 3696 0 _019_
rlabel metal3 100184 5096 100184 5096 0 _020_
rlabel metal2 101192 5936 101192 5936 0 _021_
rlabel metal2 98112 5320 98112 5320 0 _022_
rlabel metal3 99344 12152 99344 12152 0 _023_
rlabel metal3 100632 12824 100632 12824 0 _024_
rlabel metal2 102200 5488 102200 5488 0 _025_
rlabel metal2 102984 5936 102984 5936 0 _026_
rlabel metal2 103768 6328 103768 6328 0 _027_
rlabel metal2 104888 5936 104888 5936 0 _028_
rlabel metal2 107128 4984 107128 4984 0 _029_
rlabel metal3 112336 5096 112336 5096 0 _030_
rlabel metal2 110376 4200 110376 4200 0 _031_
rlabel metal2 110712 18256 110712 18256 0 _032_
rlabel metal2 112056 5320 112056 5320 0 _033_
rlabel metal2 114184 5600 114184 5600 0 _034_
rlabel metal2 117768 5432 117768 5432 0 _035_
rlabel metal2 116200 5936 116200 5936 0 _036_
rlabel metal2 119000 4928 119000 4928 0 _037_
rlabel metal3 119112 4984 119112 4984 0 _038_
rlabel metal3 119448 5880 119448 5880 0 _039_
rlabel metal3 131936 4984 131936 4984 0 _040_
rlabel metal2 125496 5432 125496 5432 0 _041_
rlabel metal2 146160 7560 146160 7560 0 addr[0]
rlabel metal3 144760 6552 144760 6552 0 addr[1]
rlabel metal2 146888 4032 146888 4032 0 addr[2]
rlabel metal3 148176 4872 148176 4872 0 addr[3]
rlabel metal2 147336 5712 147336 5712 0 addr[4]
rlabel metal3 148106 6552 148106 6552 0 addr[5]
rlabel metal2 147000 7728 147000 7728 0 addr[6]
rlabel metal3 148050 8344 148050 8344 0 addr[7]
rlabel metal2 147000 9408 147000 9408 0 addr[8]
rlabel metal2 146888 10304 146888 10304 0 addr[9]
rlabel metal2 6888 854 6888 854 0 addr_mem0[0]
rlabel metal2 8568 2198 8568 2198 0 addr_mem0[1]
rlabel metal2 10248 2198 10248 2198 0 addr_mem0[2]
rlabel metal2 11928 2198 11928 2198 0 addr_mem0[3]
rlabel metal2 13608 2086 13608 2086 0 addr_mem0[4]
rlabel metal2 15288 2086 15288 2086 0 addr_mem0[5]
rlabel metal2 16968 854 16968 854 0 addr_mem0[6]
rlabel metal2 18648 2478 18648 2478 0 addr_mem0[7]
rlabel metal2 20328 2198 20328 2198 0 addr_mem0[8]
rlabel metal2 77448 2198 77448 2198 0 addr_mem1[0]
rlabel metal2 79128 2198 79128 2198 0 addr_mem1[1]
rlabel metal2 80808 2366 80808 2366 0 addr_mem1[2]
rlabel metal2 82488 2086 82488 2086 0 addr_mem1[3]
rlabel metal2 84168 2086 84168 2086 0 addr_mem1[4]
rlabel metal3 86296 3864 86296 3864 0 addr_mem1[5]
rlabel metal3 88144 3640 88144 3640 0 addr_mem1[6]
rlabel metal3 89880 3640 89880 3640 0 addr_mem1[7]
rlabel metal3 91336 4200 91336 4200 0 addr_mem1[8]
rlabel metal3 146440 5768 146440 5768 0 csb
rlabel metal2 5208 2086 5208 2086 0 csb_mem0
rlabel metal2 75768 2198 75768 2198 0 csb_mem1
rlabel metal2 146104 11200 146104 11200 0 dout[0]
rlabel metal3 147658 19992 147658 19992 0 dout[10]
rlabel metal2 146104 21168 146104 21168 0 dout[11]
rlabel metal2 146104 22008 146104 22008 0 dout[12]
rlabel metal2 146104 22848 146104 22848 0 dout[13]
rlabel metal2 146104 23744 146104 23744 0 dout[14]
rlabel metal2 146104 24528 146104 24528 0 dout[15]
rlabel metal3 147658 25368 147658 25368 0 dout[16]
rlabel metal2 146104 26600 146104 26600 0 dout[17]
rlabel metal2 146104 27440 146104 27440 0 dout[18]
rlabel metal2 146104 28336 146104 28336 0 dout[19]
rlabel metal2 146104 11984 146104 11984 0 dout[1]
rlabel metal2 146104 29120 146104 29120 0 dout[20]
rlabel metal2 146104 30016 146104 30016 0 dout[21]
rlabel metal2 146104 30800 146104 30800 0 dout[22]
rlabel metal3 147658 31640 147658 31640 0 dout[23]
rlabel metal2 146104 32872 146104 32872 0 dout[24]
rlabel metal2 146104 33712 146104 33712 0 dout[25]
rlabel metal2 146104 34552 146104 34552 0 dout[26]
rlabel metal2 146104 35392 146104 35392 0 dout[27]
rlabel metal2 145992 36288 145992 36288 0 dout[28]
rlabel metal2 147784 36792 147784 36792 0 dout[29]
rlabel metal3 147658 12824 147658 12824 0 dout[2]
rlabel metal2 144368 36568 144368 36568 0 dout[30]
rlabel metal2 147672 37184 147672 37184 0 dout[31]
rlabel metal2 146104 14056 146104 14056 0 dout[3]
rlabel metal2 146104 14896 146104 14896 0 dout[4]
rlabel metal2 146104 15736 146104 15736 0 dout[5]
rlabel metal2 146104 16632 146104 16632 0 dout[6]
rlabel metal2 146104 17472 146104 17472 0 dout[7]
rlabel metal2 146104 18256 146104 18256 0 dout[8]
rlabel metal3 147658 19096 147658 19096 0 dout[9]
rlabel metal2 21896 4200 21896 4200 0 dout_mem0[0]
rlabel metal2 38864 3416 38864 3416 0 dout_mem0[10]
rlabel metal2 40656 4200 40656 4200 0 dout_mem0[11]
rlabel metal2 42056 3416 42056 3416 0 dout_mem0[12]
rlabel metal2 43848 2590 43848 2590 0 dout_mem0[13]
rlabel metal2 45696 4424 45696 4424 0 dout_mem0[14]
rlabel metal2 47096 3416 47096 3416 0 dout_mem0[15]
rlabel metal2 48888 2478 48888 2478 0 dout_mem0[16]
rlabel metal2 50624 3416 50624 3416 0 dout_mem0[17]
rlabel metal2 52136 4200 52136 4200 0 dout_mem0[18]
rlabel metal2 53816 3416 53816 3416 0 dout_mem0[19]
rlabel metal2 23576 3416 23576 3416 0 dout_mem0[1]
rlabel metal2 55608 2590 55608 2590 0 dout_mem0[20]
rlabel metal2 57288 2086 57288 2086 0 dout_mem0[21]
rlabel metal2 58856 3416 58856 3416 0 dout_mem0[22]
rlabel metal2 60536 4200 60536 4200 0 dout_mem0[23]
rlabel metal2 62384 3416 62384 3416 0 dout_mem0[24]
rlabel metal2 63784 4984 63784 4984 0 dout_mem0[25]
rlabel metal2 65576 3416 65576 3416 0 dout_mem0[26]
rlabel metal2 67368 2590 67368 2590 0 dout_mem0[27]
rlabel metal2 69216 4424 69216 4424 0 dout_mem0[28]
rlabel metal2 70672 3416 70672 3416 0 dout_mem0[29]
rlabel metal2 25200 4200 25200 4200 0 dout_mem0[2]
rlabel metal2 72520 4200 72520 4200 0 dout_mem0[30]
rlabel metal2 74536 4592 74536 4592 0 dout_mem0[31]
rlabel metal2 27104 3416 27104 3416 0 dout_mem0[3]
rlabel metal2 28728 2590 28728 2590 0 dout_mem0[4]
rlabel metal2 30576 4424 30576 4424 0 dout_mem0[5]
rlabel metal2 32088 2086 32088 2086 0 dout_mem0[6]
rlabel metal2 33936 4424 33936 4424 0 dout_mem0[7]
rlabel metal2 35336 3416 35336 3416 0 dout_mem0[8]
rlabel metal2 37016 4200 37016 4200 0 dout_mem0[9]
rlabel metal2 92736 3416 92736 3416 0 dout_mem1[0]
rlabel metal2 110936 4032 110936 4032 0 dout_mem1[10]
rlabel metal2 112616 3472 112616 3472 0 dout_mem1[11]
rlabel metal3 113344 3416 113344 3416 0 dout_mem1[12]
rlabel metal2 114856 2800 114856 2800 0 dout_mem1[13]
rlabel metal2 116256 4424 116256 4424 0 dout_mem1[14]
rlabel metal3 118160 3416 118160 3416 0 dout_mem1[15]
rlabel metal3 120064 3416 120064 3416 0 dout_mem1[16]
rlabel metal3 121576 3416 121576 3416 0 dout_mem1[17]
rlabel metal2 122752 3416 122752 3416 0 dout_mem1[18]
rlabel metal2 124376 4200 124376 4200 0 dout_mem1[19]
rlabel metal3 94304 4424 94304 4424 0 dout_mem1[1]
rlabel metal2 126112 3416 126112 3416 0 dout_mem1[20]
rlabel metal2 127848 3262 127848 3262 0 dout_mem1[21]
rlabel metal2 132216 3472 132216 3472 0 dout_mem1[22]
rlabel metal2 132440 3920 132440 3920 0 dout_mem1[23]
rlabel metal3 133672 4424 133672 4424 0 dout_mem1[24]
rlabel metal3 135352 3416 135352 3416 0 dout_mem1[25]
rlabel metal2 138040 3920 138040 3920 0 dout_mem1[26]
rlabel metal3 138600 4200 138600 4200 0 dout_mem1[27]
rlabel metal3 140280 3416 140280 3416 0 dout_mem1[28]
rlabel metal3 141568 3416 141568 3416 0 dout_mem1[29]
rlabel metal3 95760 3416 95760 3416 0 dout_mem1[2]
rlabel metal3 143584 3416 143584 3416 0 dout_mem1[30]
rlabel metal2 144480 4984 144480 4984 0 dout_mem1[31]
rlabel metal3 97832 3416 97832 3416 0 dout_mem1[3]
rlabel metal2 99232 3416 99232 3416 0 dout_mem1[4]
rlabel metal2 100856 4200 100856 4200 0 dout_mem1[5]
rlabel metal2 103096 2800 103096 2800 0 dout_mem1[6]
rlabel metal3 105560 3528 105560 3528 0 dout_mem1[7]
rlabel metal3 107352 3416 107352 3416 0 dout_mem1[8]
rlabel metal2 108024 3752 108024 3752 0 dout_mem1[9]
rlabel metal2 77672 5320 77672 5320 0 net1
rlabel metal2 145208 9016 145208 9016 0 net10
rlabel metal3 141904 23016 141904 23016 0 net100
rlabel metal2 119336 5992 119336 5992 0 net101
rlabel metal2 120232 5880 120232 5880 0 net102
rlabel metal3 121184 25144 121184 25144 0 net103
rlabel metal2 144984 26992 144984 26992 0 net104
rlabel metal2 144984 27776 144984 27776 0 net105
rlabel metal3 142744 28616 142744 28616 0 net106
rlabel metal2 101528 7112 101528 7112 0 net107
rlabel metal2 144984 29344 144984 29344 0 net108
rlabel metal3 141512 29960 141512 29960 0 net109
rlabel metal2 76216 6608 76216 6608 0 net11
rlabel metal2 144984 30912 144984 30912 0 net110
rlabel metal2 144984 31640 144984 31640 0 net111
rlabel metal2 144984 33208 144984 33208 0 net112
rlabel metal2 144984 34048 144984 34048 0 net113
rlabel metal3 142856 34664 142856 34664 0 net114
rlabel metal3 143248 35560 143248 35560 0 net115
rlabel metal2 144032 35560 144032 35560 0 net116
rlabel metal3 143528 7672 143528 7672 0 net117
rlabel metal2 144424 12264 144424 12264 0 net118
rlabel metal3 140616 36232 140616 36232 0 net119
rlabel metal2 23744 4200 23744 4200 0 net12
rlabel metal3 143080 3304 143080 3304 0 net120
rlabel metal2 100520 13328 100520 13328 0 net121
rlabel metal2 144312 14000 144312 14000 0 net122
rlabel metal2 144984 15960 144984 15960 0 net123
rlabel metal3 144648 16856 144648 16856 0 net124
rlabel metal2 144984 17528 144984 17528 0 net125
rlabel metal2 115864 16688 115864 16688 0 net126
rlabel metal3 144200 18984 144200 18984 0 net127
rlabel metal2 40320 3640 40320 3640 0 net13
rlabel metal2 43064 3528 43064 3528 0 net14
rlabel metal2 43736 2352 43736 2352 0 net15
rlabel metal2 45192 2856 45192 2856 0 net16
rlabel metal3 115696 5992 115696 5992 0 net17
rlabel metal2 48104 3192 48104 3192 0 net18
rlabel metal2 51016 5880 51016 5880 0 net19
rlabel metal2 78904 4760 78904 4760 0 net2
rlabel metal2 52080 3640 52080 3640 0 net20
rlabel metal3 122528 5992 122528 5992 0 net21
rlabel metal2 124936 3976 124936 3976 0 net22
rlabel metal2 24584 2632 24584 2632 0 net23
rlabel metal2 56896 4200 56896 4200 0 net24
rlabel metal2 59024 4200 59024 4200 0 net25
rlabel metal2 59864 5264 59864 5264 0 net26
rlabel metal2 62216 3360 62216 3360 0 net27
rlabel metal2 63840 3640 63840 3640 0 net28
rlabel metal2 134008 6048 134008 6048 0 net29
rlabel metal2 142072 3416 142072 3416 0 net3
rlabel metal2 67256 2296 67256 2296 0 net30
rlabel metal2 68712 2800 68712 2800 0 net31
rlabel metal2 70616 5096 70616 5096 0 net32
rlabel metal2 140000 6664 140000 6664 0 net33
rlabel metal2 27160 4760 27160 4760 0 net34
rlabel metal2 74760 7336 74760 7336 0 net35
rlabel metal2 75600 3640 75600 3640 0 net36
rlabel metal2 28560 3640 28560 3640 0 net37
rlabel metal2 30072 5040 30072 5040 0 net38
rlabel metal2 101864 3640 101864 3640 0 net39
rlabel metal2 144816 5208 144816 5208 0 net4
rlabel metal2 101976 6048 101976 6048 0 net40
rlabel metal2 35560 4200 35560 4200 0 net41
rlabel metal2 36344 5432 36344 5432 0 net42
rlabel metal2 38696 3416 38696 3416 0 net43
rlabel metal2 105672 5432 105672 5432 0 net44
rlabel metal2 110152 4928 110152 4928 0 net45
rlabel metal2 111944 3640 111944 3640 0 net46
rlabel metal2 113848 4648 113848 4648 0 net47
rlabel metal2 115864 4368 115864 4368 0 net48
rlabel metal2 116760 4928 116760 4928 0 net49
rlabel metal2 144984 5992 144984 5992 0 net5
rlabel metal2 117992 4648 117992 4648 0 net50
rlabel metal2 118776 4648 118776 4648 0 net51
rlabel metal2 122808 4648 122808 4648 0 net52
rlabel metal2 123592 4648 123592 4648 0 net53
rlabel metal2 125944 4648 125944 4648 0 net54
rlabel metal2 95928 4648 95928 4648 0 net55
rlabel metal3 128072 4088 128072 4088 0 net56
rlabel metal2 129416 4648 129416 4648 0 net57
rlabel metal2 130368 5656 130368 5656 0 net58
rlabel metal2 131432 4648 131432 4648 0 net59
rlabel metal2 122696 6944 122696 6944 0 net6
rlabel metal2 132328 4928 132328 4928 0 net60
rlabel metal2 135128 4368 135128 4368 0 net61
rlabel metal2 137032 4648 137032 4648 0 net62
rlabel metal2 138936 4368 138936 4368 0 net63
rlabel metal2 141456 4200 141456 4200 0 net64
rlabel metal2 140840 4928 140840 4928 0 net65
rlabel metal2 97720 3640 97720 3640 0 net66
rlabel metal2 138936 6664 138936 6664 0 net67
rlabel metal3 140952 5656 140952 5656 0 net68
rlabel metal2 98224 5656 98224 5656 0 net69
rlabel metal2 144760 7280 144760 7280 0 net7
rlabel metal2 99792 5096 99792 5096 0 net70
rlabel metal2 102648 4648 102648 4648 0 net71
rlabel metal2 103432 4648 103432 4648 0 net72
rlabel metal2 104552 4648 104552 4648 0 net73
rlabel metal2 106456 4368 106456 4368 0 net74
rlabel metal2 109704 4200 109704 4200 0 net75
rlabel metal3 74760 4424 74760 4424 0 net76
rlabel metal2 78008 5936 78008 5936 0 net77
rlabel metal3 11760 4536 11760 4536 0 net78
rlabel metal3 14056 4536 14056 4536 0 net79
rlabel metal2 90328 7056 90328 7056 0 net8
rlabel metal2 14952 3640 14952 3640 0 net80
rlabel metal2 16912 3528 16912 3528 0 net81
rlabel metal3 73080 3584 73080 3584 0 net82
rlabel metal2 20552 4144 20552 4144 0 net83
rlabel metal2 21448 3752 21448 3752 0 net84
rlabel metal2 77504 4424 77504 4424 0 net85
rlabel metal2 79240 3976 79240 3976 0 net86
rlabel metal2 81704 3976 81704 3976 0 net87
rlabel metal2 82488 4592 82488 4592 0 net88
rlabel metal2 84840 3976 84840 3976 0 net89
rlabel metal2 90776 7560 90776 7560 0 net9
rlabel metal2 85848 4592 85848 4592 0 net90
rlabel metal2 88200 3976 88200 3976 0 net91
rlabel metal2 89656 3976 89656 3976 0 net92
rlabel metal3 90832 4424 90832 4424 0 net93
rlabel metal2 7000 3416 7000 3416 0 net94
rlabel metal2 75824 4872 75824 4872 0 net95
rlabel metal2 144424 10976 144424 10976 0 net96
rlabel metal2 144984 20664 144984 20664 0 net97
rlabel metal3 123144 5880 123144 5880 0 net98
rlabel metal2 144984 22232 144984 22232 0 net99
<< properties >>
string FIXED_BBOX 0 0 150000 40000
<< end >>
