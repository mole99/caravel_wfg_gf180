// This is the unpowered netlist.
module merge_memory (csb,
    csb_mem0,
    csb_mem1,
    addr,
    addr_mem0,
    addr_mem1,
    dout,
    dout_mem0,
    dout_mem1);
 input csb;
 output csb_mem0;
 output csb_mem1;
 input [9:0] addr;
 output [8:0] addr_mem0;
 output [8:0] addr_mem1;
 output [31:0] dout;
 input [31:0] dout_mem0;
 input [31:0] dout_mem1;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _042_ (.I(net10),
    .Z(_040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _043_ (.I(_040_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _044_ (.I0(net20),
    .I1(net52),
    .S(_041_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _045_ (.I(_000_),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _046_ (.I0(net21),
    .I1(net53),
    .S(_041_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _047_ (.I(_001_),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _048_ (.I0(net22),
    .I1(net54),
    .S(_041_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _049_ (.I(_002_),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _050_ (.I0(net24),
    .I1(net56),
    .S(_041_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _051_ (.I(_003_),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _052_ (.I(_040_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _053_ (.I0(net25),
    .I1(net57),
    .S(_004_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _054_ (.I(_005_),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _055_ (.I0(net26),
    .I1(net58),
    .S(_004_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _056_ (.I(_006_),
    .Z(net110));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _057_ (.I0(net27),
    .I1(net59),
    .S(_004_),
    .Z(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _058_ (.I(_007_),
    .Z(net111));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _059_ (.I0(net28),
    .I1(net60),
    .S(_004_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _060_ (.I(_008_),
    .Z(net112));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _061_ (.I(_040_),
    .Z(_009_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _062_ (.I0(net29),
    .I1(net61),
    .S(_009_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _063_ (.I(_010_),
    .Z(net113));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _064_ (.I0(net30),
    .I1(net62),
    .S(_009_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _065_ (.I(_011_),
    .Z(net114));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _066_ (.I0(net31),
    .I1(net63),
    .S(_009_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _067_ (.I(_012_),
    .Z(net115));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _068_ (.I0(net32),
    .I1(net64),
    .S(_009_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _069_ (.I(_013_),
    .Z(net116));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _070_ (.I(_040_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _071_ (.I0(net33),
    .I1(net65),
    .S(_014_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _072_ (.I(_015_),
    .Z(net117));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _073_ (.I0(net35),
    .I1(net67),
    .S(_014_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _074_ (.I(_016_),
    .Z(net119));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _075_ (.I0(net36),
    .I1(net68),
    .S(_014_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _076_ (.I(_017_),
    .Z(net120));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _077_ (.I0(net12),
    .I1(net44),
    .S(_014_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _078_ (.I(_018_),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _079_ (.I(net10),
    .Z(_019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _080_ (.I(_019_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _081_ (.I0(net23),
    .I1(net55),
    .S(_020_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _082_ (.I(_021_),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _083_ (.I0(net34),
    .I1(net66),
    .S(_020_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _084_ (.I(_022_),
    .Z(net118));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _085_ (.I0(net37),
    .I1(net69),
    .S(_020_),
    .Z(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _086_ (.I(_023_),
    .Z(net121));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _087_ (.I0(net38),
    .I1(net70),
    .S(_020_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _088_ (.I(_024_),
    .Z(net122));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _089_ (.I(_019_),
    .Z(_025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _090_ (.I0(net39),
    .I1(net71),
    .S(_025_),
    .Z(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _091_ (.I(_026_),
    .Z(net123));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _092_ (.I0(net40),
    .I1(net72),
    .S(_025_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _093_ (.I(_027_),
    .Z(net124));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _094_ (.I0(net41),
    .I1(net73),
    .S(_025_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _095_ (.I(_028_),
    .Z(net125));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _096_ (.I0(net42),
    .I1(net74),
    .S(_025_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _097_ (.I(_029_),
    .Z(net126));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _098_ (.I(_019_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _099_ (.I0(net43),
    .I1(net75),
    .S(_030_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _100_ (.I(_031_),
    .Z(net127));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _101_ (.I0(net13),
    .I1(net45),
    .S(_030_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _102_ (.I(_032_),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _103_ (.I0(net14),
    .I1(net46),
    .S(_030_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _104_ (.I(_033_),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _105_ (.I0(net15),
    .I1(net47),
    .S(_030_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _106_ (.I(_034_),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _107_ (.I(_019_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _108_ (.I0(net16),
    .I1(net48),
    .S(_035_),
    .Z(_036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _109_ (.I(_036_),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _110_ (.I0(net17),
    .I1(net49),
    .S(_035_),
    .Z(_037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _111_ (.I(_037_),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _112_ (.I0(net18),
    .I1(net50),
    .S(_035_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _113_ (.I(_038_),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _114_ (.I0(net19),
    .I1(net51),
    .S(_035_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _115_ (.I(_039_),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _116_ (.I(net1),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _117_ (.I(net2),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _118_ (.I(net3),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _119_ (.I(net4),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _120_ (.I(net5),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _121_ (.I(net6),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _122_ (.I(net7),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _123_ (.I(net8),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _124_ (.I(net9),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _125_ (.I(net1),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _126_ (.I(net2),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _127_ (.I(net3),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _128_ (.I(net4),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _129_ (.I(net5),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _130_ (.I(net6),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _131_ (.I(net7),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _132_ (.I(net8),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _133_ (.I(net9),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _134_ (.I(net11),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _135_ (.I(net11),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_86 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_87 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_88 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_89 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_90 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_91 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_92 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_93 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_94 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_95 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_96 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_97 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_98 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(addr[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(addr[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(addr[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(addr[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(addr[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(addr[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(addr[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(addr[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(addr[8]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(addr[9]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input11 (.I(csb),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(dout_mem0[0]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input13 (.I(dout_mem0[10]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input14 (.I(dout_mem0[11]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(dout_mem0[12]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(dout_mem0[13]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(dout_mem0[14]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(dout_mem0[15]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(dout_mem0[16]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(dout_mem0[17]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(dout_mem0[18]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(dout_mem0[19]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(dout_mem0[1]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(dout_mem0[20]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(dout_mem0[21]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(dout_mem0[22]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(dout_mem0[23]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(dout_mem0[24]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(dout_mem0[25]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(dout_mem0[26]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(dout_mem0[27]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(dout_mem0[28]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(dout_mem0[29]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(dout_mem0[2]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(dout_mem0[30]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(dout_mem0[31]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(dout_mem0[3]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(dout_mem0[4]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input39 (.I(dout_mem0[5]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(dout_mem0[6]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(dout_mem0[7]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(dout_mem0[8]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(dout_mem0[9]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input44 (.I(dout_mem1[0]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input45 (.I(dout_mem1[10]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input46 (.I(dout_mem1[11]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input47 (.I(dout_mem1[12]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input48 (.I(dout_mem1[13]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input49 (.I(dout_mem1[14]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input50 (.I(dout_mem1[15]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input51 (.I(dout_mem1[16]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input52 (.I(dout_mem1[17]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input53 (.I(dout_mem1[18]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input54 (.I(dout_mem1[19]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input55 (.I(dout_mem1[1]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input56 (.I(dout_mem1[20]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input57 (.I(dout_mem1[21]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input58 (.I(dout_mem1[22]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input59 (.I(dout_mem1[23]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input60 (.I(dout_mem1[24]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input61 (.I(dout_mem1[25]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input62 (.I(dout_mem1[26]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input63 (.I(dout_mem1[27]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input64 (.I(dout_mem1[28]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input65 (.I(dout_mem1[29]),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input66 (.I(dout_mem1[2]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input67 (.I(dout_mem1[30]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input68 (.I(dout_mem1[31]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input69 (.I(dout_mem1[3]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input70 (.I(dout_mem1[4]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input71 (.I(dout_mem1[5]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input72 (.I(dout_mem1[6]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input73 (.I(dout_mem1[7]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input74 (.I(dout_mem1[8]),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input75 (.I(dout_mem1[9]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output76 (.I(net76),
    .Z(addr_mem0[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output77 (.I(net77),
    .Z(addr_mem0[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output78 (.I(net78),
    .Z(addr_mem0[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output79 (.I(net79),
    .Z(addr_mem0[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output80 (.I(net80),
    .Z(addr_mem0[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output81 (.I(net81),
    .Z(addr_mem0[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output82 (.I(net82),
    .Z(addr_mem0[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output83 (.I(net83),
    .Z(addr_mem0[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output84 (.I(net84),
    .Z(addr_mem0[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output85 (.I(net85),
    .Z(addr_mem1[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output86 (.I(net86),
    .Z(addr_mem1[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output87 (.I(net87),
    .Z(addr_mem1[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output88 (.I(net88),
    .Z(addr_mem1[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output89 (.I(net89),
    .Z(addr_mem1[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output90 (.I(net90),
    .Z(addr_mem1[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output91 (.I(net91),
    .Z(addr_mem1[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output92 (.I(net92),
    .Z(addr_mem1[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output93 (.I(net93),
    .Z(addr_mem1[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output94 (.I(net94),
    .Z(csb_mem0));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output95 (.I(net95),
    .Z(csb_mem1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output96 (.I(net96),
    .Z(dout[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output97 (.I(net97),
    .Z(dout[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output98 (.I(net98),
    .Z(dout[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output99 (.I(net99),
    .Z(dout[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output100 (.I(net100),
    .Z(dout[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output101 (.I(net101),
    .Z(dout[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output102 (.I(net102),
    .Z(dout[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output103 (.I(net103),
    .Z(dout[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output104 (.I(net104),
    .Z(dout[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output105 (.I(net105),
    .Z(dout[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output106 (.I(net106),
    .Z(dout[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output107 (.I(net107),
    .Z(dout[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output108 (.I(net108),
    .Z(dout[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output109 (.I(net109),
    .Z(dout[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output110 (.I(net110),
    .Z(dout[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output111 (.I(net111),
    .Z(dout[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output112 (.I(net112),
    .Z(dout[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output113 (.I(net113),
    .Z(dout[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output114 (.I(net114),
    .Z(dout[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output115 (.I(net115),
    .Z(dout[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output116 (.I(net116),
    .Z(dout[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output117 (.I(net117),
    .Z(dout[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output118 (.I(net118),
    .Z(dout[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output119 (.I(net119),
    .Z(dout[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output120 (.I(net120),
    .Z(dout[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output121 (.I(net121),
    .Z(dout[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output122 (.I(net122),
    .Z(dout[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output123 (.I(net123),
    .Z(dout[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output124 (.I(net124),
    .Z(dout[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output125 (.I(net125),
    .Z(dout[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output126 (.I(net126),
    .Z(dout[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output127 (.I(net127),
    .Z(dout[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__077__S (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__075__S (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__073__S (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__071__S (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__107__I (.I(_019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__098__I (.I(_019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__089__I (.I(_019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__080__I (.I(_019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__086__I (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__102__I (.I(_032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__070__I (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__061__I (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__052__I (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__043__I (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(csb));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(dout_mem0[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(dout_mem0[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(dout_mem0[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(dout_mem0[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(dout_mem0[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(dout_mem0[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(dout_mem0[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(dout_mem0[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(dout_mem0[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(dout_mem0[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(dout_mem0[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(dout_mem0[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(dout_mem0[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(dout_mem0[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(dout_mem0[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(dout_mem0[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(dout_mem0[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(dout_mem0[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(dout_mem0[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(dout_mem0[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(dout_mem0[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(dout_mem0[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(dout_mem0[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(dout_mem0[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(dout_mem0[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(dout_mem0[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(dout_mem0[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(dout_mem0[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(dout_mem0[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(dout_mem0[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(dout_mem0[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(dout_mem0[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(dout_mem1[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(dout_mem1[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(dout_mem1[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(dout_mem1[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(dout_mem1[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(dout_mem1[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(dout_mem1[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(dout_mem1[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(dout_mem1[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(dout_mem1[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(dout_mem1[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(dout_mem1[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(dout_mem1[20]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(dout_mem1[21]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(dout_mem1[22]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(dout_mem1[23]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(dout_mem1[24]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(dout_mem1[25]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(dout_mem1[26]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(dout_mem1[27]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(dout_mem1[28]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(dout_mem1[29]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(dout_mem1[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(dout_mem1[30]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(dout_mem1[31]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(dout_mem1[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(dout_mem1[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(dout_mem1[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(dout_mem1[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(dout_mem1[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(dout_mem1[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(dout_mem1[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__125__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__116__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__126__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__117__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__127__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__118__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__128__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__119__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__129__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__120__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__130__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__121__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__131__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__122__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__132__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__123__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__133__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__124__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__079__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__042__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__135__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__134__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__077__I0 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__101__I0 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__103__I0 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__105__I0 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__108__I0 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__110__I0 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__112__I0 (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__114__I0 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__044__I0 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__046__I0 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__048__I0 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__081__I0 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__050__I0 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__053__I0 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__055__I0 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__057__I0 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__059__I0 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__062__I0 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__064__I0 (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__066__I0 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__068__I0 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__071__I0 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__083__I0 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__073__I0 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__075__I0 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__085__I0 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__087__I0 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__090__I0 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__092__I0 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__094__I0 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__096__I0 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__099__I0 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__077__I1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output76_I (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output77_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output78_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output79_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output80_I (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output81_I (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output82_I (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output83_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output84_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output94_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output96_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output100_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output101_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output102_I (.I(net102));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output103_I (.I(net103));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output104_I (.I(net104));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output105_I (.I(net105));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output106_I (.I(net106));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output107_I (.I(net107));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output108_I (.I(net108));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output109_I (.I(net109));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output110_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output111_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output112_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output113_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output114_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output115_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output116_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output117_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output118_I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output120_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output121_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output122_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output123_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output124_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output125_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output126_I (.I(net126));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output127_I (.I(net127));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
endmodule

